/*
  Eric Villasenor
  evillase@gmail.com

  this block is the coherence protocol
  and artibtration for ram
*/

// interface include
`include "control_unit_if.vh"

// memory types
`include "cpu_types_pkg.vh"

module control_unit
  (
   control_unit_if cuif
   );

   import cpu_types_pkg::*;

   r_t rtype;  //three different type of instruction
   j_t jtype;
   i_t itype;

   assign rtype = cuif.instr;
   assign jtype = cuif.instr;
   assign itype = cuif.instr;

   always_comb begin
      cuif.source1 = 0;
      cuif.source2 = 0;
      cuif.source3 = 0;
      cuif.immediate = 0;
      cuif.j_addr = 0;
      cuif.jregaddr = 0;
      cuif.aluop = ALU_ADD;
      cuif.WEN = 0;
      cuif.wdat = 0;
      cuif.wsel = 0;
      cuif.rsel1 = 0;
      cuif.rsel2 = 0;
      cuif.extop = 0;
      cuif.irsel = 0;
      cuif.memtoreg = 0;
      cuif.datamemstore = 0;
      cuif.datamemaddr = 0;
      cuif.dWEN = 0;
      cuif.dREN = 0;
      cuif.halt = 0;

      casez (itype.opcode) //I-type instruction opcode
	BEQ : begin
	   cuif.source1 = cuif.zeroflag;  //if it is zero, then branch
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.aluop = ALU_SUB;
	   cuif.WEN = 0;
	   cuif.rsel1 = itype.rs;
	   cuif.rsel2 = itype.rt;
	   cuif.irsel = 0;
	end // case: BEQ
	BNE : begin
	   cuif.source1 = ~cuif.zeroflag;  //if it is zero, then branch
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.aluop = ALU_SUB;
	   cuif.WEN = 0;
	   cuif.rsel1 = itype.rs;
	   cuif.rsel2 = itype.rt;
	   cuif.irsel = 0;  //will use rdata2 to be the second input to ALU
	end // case: BNE
	ADDI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.aluop = ALU_ADD;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.extop = 1; //will use sign extend
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	ADDIU : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 1; //will use sign extend
	   cuif.aluop = ALU_ADD;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	SLTI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 1; //will use sign extend
	   cuif.aluop = ALU_SLT;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	SLTIU : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 0; //will use UNsign extend
	   cuif.aluop = ALU_SLT;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	ANDI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 0; //will use sign extend
	   cuif.aluop = ALU_AND;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	ORI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 0; //will use sign extend
	   cuif.aluop = ALU_OR;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
   	XORI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 0; //will use sign extend
	   cuif.aluop = ALU_XOR;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
   	LUI : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 0;  //zero mean write the value of reg to mem
	   cuif.rsel1 = '0;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 2; 
	   cuif.aluop = ALU_ADD;
	   cuif.wdat = cuif.porto; //the write data into the reg from ALU output
	end // case: ADDI
	LW : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 1;  //!!!!!!!!!!!!!!!DOUBLE CHECK
	   cuif.rsel1 = itype.rs;
	   cuif.wsel = itype.rt;
	   cuif.WEN = 1;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 1; //will use sign extend
	   cuif.aluop = ALU_ADD;

	   cuif.dREN = 1;
	   cuif.datamemaddr = cuif.porto;
	end // case: ADDI
	SW : begin
	   cuif.irsel = 1;
	   cuif.memtoreg = 1; 
	   cuif.rsel1 = itype.rs;
	   cuif.rsel2 = itype.rt;
	   cuif.WEN = 0;  //will write the output into another register
	   cuif.source1 = 0;  
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = itype.imm;
	   cuif.extop = 1; //will use sign extend
	   cuif.aluop = ALU_ADD;

	   cuif.dWEN = 1;
	   cuif.datamemaddr = cuif.porto;
	   cuif.datamemstore = cuif.rdat2;
	end // case: ADDI
	HALT : begin
	   cuif.halt = 1;
	end
	J: begin
	   cuif.irsel = 0;
	   cuif.memtoreg = 0;
	   cuif.WEN = 0;
	   cuif.source1 = 0;
	   cuif.source2 = 1;
	   cuif.source3 = 0;
	   cuif.aluop = ALU_ADD;
	   cuif.j_addr = jtype.addr;
	end
	JAL: begin
	   cuif.irsel = 0;
	   cuif.memtoreg = 2;
	   cuif.WEN = 1;
	   cuif.wsel = 31; //default return register
	   cuif.source1 = 0;
	   cuif.source2 = 1;
	   cuif.source3 = 0;
	   cuif.aluop = ALU_ADD;
	   cuif.j_addr = jtype.addr;
	end // case: JAL
	RTYPE : begin
	   cuif.source1 = 0;
	   cuif.source2 = 0;
	   cuif.source3 = 0;
	   cuif.immediate = 0;
	   cuif.j_addr = 0;
	   cuif.jregaddr = 0;
	   cuif.aluop = ALU_ADD;
	   cuif.WEN = 0;
	   cuif.wdat = 0;
	   cuif.wsel = 0;
	   cuif.rsel1 = 0;
	   cuif.rsel2 = 0;
	   cuif.extop = 0;
	   cuif.irsel = 0;
	   cuif.memtoreg = 0;
	   cuif.datamemstore = 0;
	   cuif.datamemaddr = 0;
	   cuif.dWEN = 0;
	   cuif.dREN = 0;
	   cuif.halt = 0;

	   casez (rtype.funct) //I-type instruction opcode
	     ADDU : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_ADD;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     AND : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_AND;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     NOR : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_NOR;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     OR : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_OR;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     SLT : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_SLT;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     SLTU : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_SLTU;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     SLL : begin
		cuif.irsel = 1;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.extop = 0;
		cuif.immediate = rtype.shamt;
		cuif.aluop = ALU_SLL;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     SRL : begin
		cuif.irsel = 1;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.extop = 0;
		cuif.immediate = rtype.shamt;
		cuif.aluop = ALU_SRL;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     SUBU : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_SUB;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     XOR : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = rtype.rt;
		cuif.wsel = rtype.rd;
		cuif.WEN = 1;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_XOR;
		cuif.wdat = cuif.porto;
	     end // case: BEQ
	     JR : begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.rsel1 = rtype.rs;
		cuif.rsel2 = '0;
		cuif.wsel = rtype.rd;
		cuif.WEN = 0;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 1;
		cuif.aluop = ALU_ADD;
		cuif.jregaddr = cuif.porto;
	     end // case: BEQ
	     default: begin
		cuif.irsel = 0;
		cuif.memtoreg = 0;
		cuif.extop = 0;
		cuif.rsel1 = '0;
		cuif.rsel2 = '0;
		cuif.WEN = 0;
		cuif.source1 = 0;
		cuif.source2 = 0;
		cuif.source3 = 0;
		cuif.aluop = ALU_ADD;
		cuif.dWEN = 0;
		cuif.dREN = 0;
		cuif.halt = 0;
	     end // case: BEQ
	   endcase // casez (rtype.funct)
	end // case: RTYPE
      endcase // casez (itype.opcode)
   end // block: CULogic
endmodule // control_unit

	   
