// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "12/06/2016 19:17:19"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_AB10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_V4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_U1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_R6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_AF11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_AE11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_T7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_T26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_AC10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_AC17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_AG21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_AE18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_U4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_R4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_U3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_AH21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_R26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_W22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_AH11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_AG11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_T22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AD17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_T25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_AF18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_T21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_T4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_V3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|PR|Memwrite_EX~q ;
wire \CPU|DP|PR|MemToReg_EX~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~16_combout ;
wire \RAM|ramif.ramload[17]~17_combout ;
wire \RAM|ramif.ramload[18]~18_combout ;
wire \RAM|ramif.ramload[19]~19_combout ;
wire \RAM|ramif.ramload[20]~20_combout ;
wire \RAM|ramif.ramload[21]~21_combout ;
wire \RAM|ramif.ramload[22]~22_combout ;
wire \RAM|ramif.ramload[23]~23_combout ;
wire \RAM|ramif.ramload[24]~24_combout ;
wire \RAM|ramif.ramload[25]~25_combout ;
wire \RAM|ramif.ramload[26]~26_combout ;
wire \RAM|ramif.ramload[27]~27_combout ;
wire \RAM|ramif.ramload[28]~28_combout ;
wire \RAM|ramif.ramload[29]~29_combout ;
wire \RAM|ramif.ramload[30]~30_combout ;
wire \RAM|ramif.ramload[31]~31_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \ramstore~0_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.addr[1]~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|halt_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|pc ;
wire [31:0] \CPU|DP|PR|Wdata_EX ;
wire [31:0] \CPU|DP|PR|Result_EX ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.\ramif.ramaddr ({\ramaddr~59_combout ,\ramaddr~61_combout ,\ramaddr~55_combout ,\ramaddr~57_combout ,\ramaddr~51_combout ,\ramaddr~53_combout ,\ramaddr~62_combout ,\ramaddr~63_combout ,\ramaddr~45_combout ,\ramaddr~47_combout ,\ramaddr~41_combout ,\ramaddr~43_combout ,
\ramaddr~37_combout ,\ramaddr~39_combout ,\ramaddr~33_combout ,\ramaddr~35_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~1_combout ,\ramaddr~3_combout }),
	.ramaddr(\ramaddr~5_combout ),
	.ramaddr1(\ramaddr~7_combout ),
	.ramaddr2(\ramaddr~9_combout ),
	.ramaddr3(\ramaddr~11_combout ),
	.ramaddr4(\ramaddr~13_combout ),
	.ramaddr5(\ramaddr~15_combout ),
	.ramaddr6(\ramaddr~17_combout ),
	.ramaddr7(\ramaddr~19_combout ),
	.ramaddr8(\ramaddr~21_combout ),
	.ramaddr9(\ramaddr~23_combout ),
	.ramaddr10(\ramaddr~25_combout ),
	.ramaddr11(\ramaddr~27_combout ),
	.ramaddr12(\ramaddr~29_combout ),
	.ramaddr13(\ramaddr~31_combout ),
	.ramaddr14(\ramaddr~48_combout ),
	.ramaddr15(\ramaddr~49_combout ),
	.ramWEN(\ramWEN~0_combout ),
	.ramREN(\ramREN~0_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.ramaddr16(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.syiftbCTRL(\syif.tbCTRL~input_o ),
	.syifaddr_25(\syif.addr[25]~input_o ),
	.syifaddr_24(\syif.addr[24]~input_o ),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline CPU(
	.Result_EX_1(\CPU|DP|PR|Result_EX [1]),
	.pc_1(\CPU|DP|pc [1]),
	.Memwrite_EX(\CPU|DP|PR|Memwrite_EX~q ),
	.MemToReg_EX(\CPU|DP|PR|MemToReg_EX~q ),
	.Result_EX_0(\CPU|DP|PR|Result_EX [0]),
	.pc_0(\CPU|DP|pc [0]),
	.Result_EX_3(\CPU|DP|PR|Result_EX [3]),
	.pc_3(\CPU|DP|pc [3]),
	.Result_EX_2(\CPU|DP|PR|Result_EX [2]),
	.pc_2(\CPU|DP|pc [2]),
	.Result_EX_5(\CPU|DP|PR|Result_EX [5]),
	.pc_5(\CPU|DP|pc [5]),
	.Result_EX_4(\CPU|DP|PR|Result_EX [4]),
	.pc_4(\CPU|DP|pc [4]),
	.Result_EX_7(\CPU|DP|PR|Result_EX [7]),
	.pc_7(\CPU|DP|pc [7]),
	.Result_EX_6(\CPU|DP|PR|Result_EX [6]),
	.pc_6(\CPU|DP|pc [6]),
	.Result_EX_9(\CPU|DP|PR|Result_EX [9]),
	.pc_9(\CPU|DP|pc [9]),
	.Result_EX_8(\CPU|DP|PR|Result_EX [8]),
	.pc_8(\CPU|DP|pc [8]),
	.Result_EX_11(\CPU|DP|PR|Result_EX [11]),
	.pc_11(\CPU|DP|pc [11]),
	.Result_EX_10(\CPU|DP|PR|Result_EX [10]),
	.pc_10(\CPU|DP|pc [10]),
	.Result_EX_13(\CPU|DP|PR|Result_EX [13]),
	.pc_13(\CPU|DP|pc [13]),
	.Result_EX_12(\CPU|DP|PR|Result_EX [12]),
	.pc_12(\CPU|DP|pc [12]),
	.Result_EX_15(\CPU|DP|PR|Result_EX [15]),
	.pc_15(\CPU|DP|pc [15]),
	.Result_EX_14(\CPU|DP|PR|Result_EX [14]),
	.pc_14(\CPU|DP|pc [14]),
	.Result_EX_17(\CPU|DP|PR|Result_EX [17]),
	.pc_17(\CPU|DP|pc [17]),
	.Result_EX_16(\CPU|DP|PR|Result_EX [16]),
	.pc_16(\CPU|DP|pc [16]),
	.Result_EX_19(\CPU|DP|PR|Result_EX [19]),
	.pc_19(\CPU|DP|pc [19]),
	.Result_EX_18(\CPU|DP|PR|Result_EX [18]),
	.pc_18(\CPU|DP|pc [18]),
	.Result_EX_21(\CPU|DP|PR|Result_EX [21]),
	.pc_21(\CPU|DP|pc [21]),
	.Result_EX_20(\CPU|DP|PR|Result_EX [20]),
	.pc_20(\CPU|DP|pc [20]),
	.Result_EX_23(\CPU|DP|PR|Result_EX [23]),
	.pc_23(\CPU|DP|pc [23]),
	.Result_EX_22(\CPU|DP|PR|Result_EX [22]),
	.pc_22(\CPU|DP|pc [22]),
	.Result_EX_25(\CPU|DP|PR|Result_EX [25]),
	.pc_25(\CPU|DP|pc [25]),
	.Result_EX_24(\CPU|DP|PR|Result_EX [24]),
	.pc_24(\CPU|DP|pc [24]),
	.Result_EX_27(\CPU|DP|PR|Result_EX [27]),
	.pc_27(\CPU|DP|pc [27]),
	.Result_EX_26(\CPU|DP|PR|Result_EX [26]),
	.pc_26(\CPU|DP|pc [26]),
	.Result_EX_29(\CPU|DP|PR|Result_EX [29]),
	.pc_29(\CPU|DP|pc [29]),
	.Result_EX_28(\CPU|DP|PR|Result_EX [28]),
	.pc_28(\CPU|DP|pc [28]),
	.Result_EX_31(\CPU|DP|PR|Result_EX [31]),
	.pc_31(\CPU|DP|pc [31]),
	.Result_EX_30(\CPU|DP|PR|Result_EX [30]),
	.pc_30(\CPU|DP|pc [30]),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.Wdata_EX_0(\CPU|DP|PR|Wdata_EX [0]),
	.Wdata_EX_1(\CPU|DP|PR|Wdata_EX [1]),
	.Wdata_EX_2(\CPU|DP|PR|Wdata_EX [2]),
	.Wdata_EX_3(\CPU|DP|PR|Wdata_EX [3]),
	.Wdata_EX_4(\CPU|DP|PR|Wdata_EX [4]),
	.Wdata_EX_5(\CPU|DP|PR|Wdata_EX [5]),
	.Wdata_EX_6(\CPU|DP|PR|Wdata_EX [6]),
	.Wdata_EX_7(\CPU|DP|PR|Wdata_EX [7]),
	.Wdata_EX_8(\CPU|DP|PR|Wdata_EX [8]),
	.Wdata_EX_9(\CPU|DP|PR|Wdata_EX [9]),
	.Wdata_EX_10(\CPU|DP|PR|Wdata_EX [10]),
	.Wdata_EX_11(\CPU|DP|PR|Wdata_EX [11]),
	.Wdata_EX_12(\CPU|DP|PR|Wdata_EX [12]),
	.Wdata_EX_13(\CPU|DP|PR|Wdata_EX [13]),
	.Wdata_EX_14(\CPU|DP|PR|Wdata_EX [14]),
	.Wdata_EX_15(\CPU|DP|PR|Wdata_EX [15]),
	.Wdata_EX_16(\CPU|DP|PR|Wdata_EX [16]),
	.Wdata_EX_17(\CPU|DP|PR|Wdata_EX [17]),
	.Wdata_EX_18(\CPU|DP|PR|Wdata_EX [18]),
	.Wdata_EX_19(\CPU|DP|PR|Wdata_EX [19]),
	.Wdata_EX_20(\CPU|DP|PR|Wdata_EX [20]),
	.Wdata_EX_21(\CPU|DP|PR|Wdata_EX [21]),
	.Wdata_EX_22(\CPU|DP|PR|Wdata_EX [22]),
	.Wdata_EX_23(\CPU|DP|PR|Wdata_EX [23]),
	.Wdata_EX_24(\CPU|DP|PR|Wdata_EX [24]),
	.Wdata_EX_25(\CPU|DP|PR|Wdata_EX [25]),
	.Wdata_EX_26(\CPU|DP|PR|Wdata_EX [26]),
	.Wdata_EX_27(\CPU|DP|PR|Wdata_EX [27]),
	.Wdata_EX_28(\CPU|DP|PR|Wdata_EX [28]),
	.Wdata_EX_29(\CPU|DP|PR|Wdata_EX [29]),
	.Wdata_EX_30(\CPU|DP|PR|Wdata_EX [30]),
	.Wdata_EX_31(\CPU|DP|PR|Wdata_EX [31]),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST(\nRST~inputclkctrl_outclk ),
	.halt_reg(\CPU|DP|halt_reg~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (Memwrite_EX1 & (((Result_EX_1)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_1))) # (!MemToReg_EX1 & (pc_1))))

	.dataa(\CPU|DP|pc [1]),
	.datab(\CPU|DP|PR|Result_EX [1]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hCCCA;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[1]~input_o ),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hF5A0;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (Memwrite_EX1 & (Result_EX_0)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_0)) # (!MemToReg_EX1 & ((pc_0)))))

	.dataa(\CPU|DP|PR|Result_EX [0]),
	.datab(\CPU|DP|pc [0]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hAAAC;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[0]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hDD88;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (MemToReg_EX1 & (Result_EX_3)) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_3)) # (!Memwrite_EX1 & ((pc_3)))))

	.dataa(\CPU|DP|PR|Result_EX [3]),
	.datab(\CPU|DP|pc [3]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hAAAC;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout )))

	.dataa(\syif.addr[3]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~4_combout ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hAFA0;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (MemToReg_EX1 & (((Result_EX_2)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_2))) # (!Memwrite_EX1 & (pc_2))))

	.dataa(\CPU|DP|pc [2]),
	.datab(\CPU|DP|PR|MemToReg_EX~q ),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|Result_EX [2]),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hFE02;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(\syif.addr[2]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hAFA0;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (Memwrite_EX1 & (((Result_EX_5)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_5))) # (!MemToReg_EX1 & (pc_5))))

	.dataa(\CPU|DP|PR|Memwrite_EX~q ),
	.datab(\CPU|DP|pc [5]),
	.datac(\CPU|DP|PR|Result_EX [5]),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hF0E4;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.addr[5]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hB8B8;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (Memwrite_EX1 & (((Result_EX_4)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_4))) # (!MemToReg_EX1 & (pc_4))))

	.dataa(\CPU|DP|PR|Memwrite_EX~q ),
	.datab(\CPU|DP|pc [4]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Result_EX [4]),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hFE04;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(\syif.addr[4]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hBB88;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (Memwrite_EX1 & (((Result_EX_7)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_7))) # (!MemToReg_EX1 & (pc_7))))

	.dataa(\CPU|DP|PR|Memwrite_EX~q ),
	.datab(\CPU|DP|pc [7]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Result_EX [7]),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hFE04;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[7]~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hF3C0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (MemToReg_EX1 & (((Result_EX_6)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_6))) # (!Memwrite_EX1 & (pc_6))))

	.dataa(\CPU|DP|pc [6]),
	.datab(\CPU|DP|PR|MemToReg_EX~q ),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|Result_EX [6]),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hFE02;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[6]~input_o ),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hF3C0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (MemToReg_EX1 & (((Result_EX_9)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_9))) # (!Memwrite_EX1 & (pc_9))))

	.dataa(\CPU|DP|pc [9]),
	.datab(\CPU|DP|PR|Result_EX [9]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hCCCA;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hF5A0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (MemToReg_EX1 & (Result_EX_8)) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_8)) # (!Memwrite_EX1 & ((pc_8)))))

	.dataa(\CPU|DP|PR|Result_EX [8]),
	.datab(\CPU|DP|pc [8]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hAAAC;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout )))

	.dataa(\syif.addr[8]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hAFA0;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (Memwrite_EX1 & (Result_EX_11)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_11)) # (!MemToReg_EX1 & ((pc_11)))))

	.dataa(\CPU|DP|PR|Result_EX [11]),
	.datab(\CPU|DP|pc [11]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hAAAC;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hF3C0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (Memwrite_EX1 & (Result_EX_10)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_10)) # (!MemToReg_EX1 & ((pc_10)))))

	.dataa(\CPU|DP|PR|Result_EX [10]),
	.datab(\CPU|DP|pc [10]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hAAAC;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(\syif.addr[10]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hBB88;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N18
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (Memwrite_EX1 & (Result_EX_13)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_13)) # (!MemToReg_EX1 & ((pc_13)))))

	.dataa(\CPU|DP|PR|Result_EX [13]),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|pc [13]),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hAAB8;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N14
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[13]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hDD88;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N6
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (MemToReg_EX1 & (((Result_EX_12)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_12))) # (!Memwrite_EX1 & (pc_12))))

	.dataa(\CPU|DP|pc [12]),
	.datab(\CPU|DP|PR|MemToReg_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [12]),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hF0E2;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N12
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[12]~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hF5A0;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N24
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (MemToReg_EX1 & (((Result_EX_15)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_15))) # (!Memwrite_EX1 & (pc_15))))

	.dataa(\CPU|DP|pc [15]),
	.datab(\CPU|DP|PR|MemToReg_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [15]),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hF0E2;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N2
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~28_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[15]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h2277;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N30
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (Memwrite_EX1 & (((Result_EX_14)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_14))) # (!MemToReg_EX1 & (pc_14))))

	.dataa(\CPU|DP|pc [14]),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [14]),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hF0E2;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N10
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[14]~input_o ),
	.datac(\ramaddr~30_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hD8D8;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (Memwrite_EX1 & (Result_EX_17)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_17)) # (!MemToReg_EX1 & ((pc_17)))))

	.dataa(\CPU|DP|PR|Result_EX [17]),
	.datab(\CPU|DP|pc [17]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hAAAC;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout )))

	.dataa(gnd),
	.datab(\syif.addr[17]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hCFC0;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (Memwrite_EX1 & (((Result_EX_16)))) # (!Memwrite_EX1 & ((MemToReg_EX1 & ((Result_EX_16))) # (!MemToReg_EX1 & (pc_16))))

	.dataa(\CPU|DP|pc [16]),
	.datab(\CPU|DP|PR|Result_EX [16]),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(\CPU|DP|PR|MemToReg_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hCCCA;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout )))

	.dataa(\syif.addr[16]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hAFA0;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (MemToReg_EX1 & (Result_EX_19)) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_19)) # (!Memwrite_EX1 & ((pc_19)))))

	.dataa(\CPU|DP|PR|Result_EX [19]),
	.datab(\CPU|DP|pc [19]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hAAAC;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(gnd),
	.datab(\syif.addr[19]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hCFC0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (MemToReg_EX1 & (((Result_EX_18)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_18))) # (!Memwrite_EX1 & (pc_18))))

	.dataa(\CPU|DP|pc [18]),
	.datab(\CPU|DP|PR|Result_EX [18]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hCCCA;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[18]~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hF3C0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (MemToReg_EX1 & (((Result_EX_21)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_21)) # (!Memwrite_EX1 & ((pc_21)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [21]),
	.datad(\CPU|DP|pc [21]),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hF1E0;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(\syif.addr[21]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hBB88;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (MemToReg_EX1 & (((Result_EX_20)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_20)) # (!Memwrite_EX1 & ((pc_20)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [20]),
	.datad(\CPU|DP|pc [20]),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hF1E0;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(\syif.addr[20]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hB8B8;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (MemToReg_EX1 & (((Result_EX_23)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_23))) # (!Memwrite_EX1 & (pc_23))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|pc [23]),
	.datad(\CPU|DP|PR|Result_EX [23]),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hFE10;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[23]~input_o ),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hF5A0;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (MemToReg_EX1 & (((Result_EX_22)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_22))) # (!Memwrite_EX1 & (pc_22))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|pc [22]),
	.datad(\CPU|DP|PR|Result_EX [22]),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hFE10;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[22]~input_o ),
	.datad(\ramaddr~46_combout ),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hF5A0;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (MemToReg_EX1 & (Result_EX_25)) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_25)) # (!Memwrite_EX1 & ((pc_25)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Result_EX [25]),
	.datac(\CPU|DP|pc [25]),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hCCD8;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (MemToReg_EX1 & (((Result_EX_24)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_24))) # (!Memwrite_EX1 & (pc_24))))

	.dataa(\CPU|DP|pc [24]),
	.datab(\CPU|DP|PR|Result_EX [24]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hCCCA;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (MemToReg_EX1 & (((Result_EX_27)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & ((Result_EX_27))) # (!Memwrite_EX1 & (pc_27))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|pc [27]),
	.datac(\CPU|DP|PR|Result_EX [27]),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hF0E4;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[27]~input_o ),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hF3C0;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (MemToReg_EX1 & (Result_EX_26)) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_26)) # (!Memwrite_EX1 & ((pc_26)))))

	.dataa(\CPU|DP|PR|Result_EX [26]),
	.datab(\CPU|DP|pc [26]),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|PR|Memwrite_EX~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hAAAC;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(\syif.addr[26]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hBB88;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (MemToReg_EX1 & (((Result_EX_29)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_29)) # (!Memwrite_EX1 & ((pc_29)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [29]),
	.datad(\CPU|DP|pc [29]),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hF1E0;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[29]~input_o ),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hF5A0;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (MemToReg_EX1 & (((Result_EX_28)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_28)) # (!Memwrite_EX1 & ((pc_28)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [28]),
	.datad(\CPU|DP|pc [28]),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hF1E0;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[28]~input_o ),
	.datad(\ramaddr~56_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hF5A0;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (MemToReg_EX1 & (((Result_EX_31)))) # (!MemToReg_EX1 & ((Memwrite_EX1 & (Result_EX_31)) # (!Memwrite_EX1 & ((pc_31)))))

	.dataa(\CPU|DP|PR|MemToReg_EX~q ),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|Result_EX [31]),
	.datad(\CPU|DP|pc [31]),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hF1E0;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[31]~input_o ),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hF5A0;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (Memwrite_EX1 & (Result_EX_30)) # (!Memwrite_EX1 & ((MemToReg_EX1 & (Result_EX_30)) # (!MemToReg_EX1 & ((pc_30)))))

	.dataa(\CPU|DP|PR|Result_EX [30]),
	.datab(\CPU|DP|PR|Memwrite_EX~q ),
	.datac(\CPU|DP|PR|MemToReg_EX~q ),
	.datad(\CPU|DP|pc [30]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hABA8;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[30]~input_o ),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hF5A0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!Memwrite_EX1)))

	.dataa(\syif.WEN~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Memwrite_EX~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h4747;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & !\syif.REN~input_o )

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(gnd),
	.datad(\syif.REN~input_o ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h00AA;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X1_Y36_N15
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[0]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_0))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [0]),
	.datad(\syif.store[0]~input_o ),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hFC30;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[25]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~48_combout ))

	.dataa(\ramaddr~48_combout ),
	.datab(\syif.addr[25]~input_o ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hCCAA;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~49_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[24]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~49_combout ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hDD88;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\syif.tbCTRL~input_o  & (\syif.store[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_1)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[1]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [1]),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hF3C0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\syif.tbCTRL~input_o  & (\syif.store[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_2)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[2]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [2]),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hF3C0;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N16
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.tbCTRL~input_o  & (\syif.store[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_3)))

	.dataa(gnd),
	.datab(\syif.store[3]~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [3]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hCCF0;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N26
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[4]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_4))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PR|Wdata_EX [4]),
	.datac(\syif.store[4]~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hE4E4;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\syif.tbCTRL~input_o  & (\syif.store[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_5)))

	.dataa(\syif.store[5]~input_o ),
	.datab(\CPU|DP|PR|Wdata_EX [5]),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hAACC;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & (\syif.store[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_6)))

	.dataa(\syif.store[6]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [6]),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hBB88;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[7]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_7))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [7]),
	.datad(\syif.store[7]~input_o ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hFC30;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.tbCTRL~input_o  & (\syif.store[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_8)))

	.dataa(\syif.store[8]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [8]),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hBB88;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\syif.tbCTRL~input_o  & (\syif.store[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_9)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[9]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [9]),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hF3C0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.tbCTRL~input_o  & (\syif.store[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_10)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[10]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hF5A0;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.tbCTRL~input_o  & (\syif.store[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_11)))

	.dataa(gnd),
	.datab(\syif.store[11]~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [11]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hCCF0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (\syif.tbCTRL~input_o  & (\syif.store[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_12)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[12]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [12]),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hF3C0;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\syif.tbCTRL~input_o  & (\syif.store[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_13)))

	.dataa(gnd),
	.datab(\syif.store[13]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [13]),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hCFC0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\syif.tbCTRL~input_o  & (\syif.store[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_14)))

	.dataa(\syif.store[14]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [14]),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hAFA0;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.tbCTRL~input_o  & (\syif.store[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_15)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[15]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [15]),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hF3C0;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\syif.tbCTRL~input_o  & (\syif.store[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_16)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[16]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [16]),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hF3C0;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\syif.tbCTRL~input_o  & (\syif.store[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_17)))

	.dataa(\syif.store[17]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [17]),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hBB88;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (\syif.tbCTRL~input_o  & (\syif.store[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_18)))

	.dataa(\syif.store[18]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [18]),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hB8B8;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\syif.tbCTRL~input_o  & (\syif.store[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_19)))

	.dataa(\syif.store[19]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hAFA0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\syif.tbCTRL~input_o  & (\syif.store[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_20)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[20]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hF3C0;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[21]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_21))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [21]),
	.datad(\syif.store[21]~input_o ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hFC30;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & (\syif.store[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_22)))

	.dataa(\syif.store[22]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [22]),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hBB88;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.tbCTRL~input_o  & (\syif.store[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_23)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[23]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [23]),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hF3C0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\syif.tbCTRL~input_o  & (\syif.store[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_24)))

	.dataa(\syif.store[24]~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|PR|Wdata_EX [24]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hAAF0;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.tbCTRL~input_o  & (\syif.store[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_25)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[25]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [25]),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hF3C0;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\syif.tbCTRL~input_o  & (\syif.store[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_26)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[26]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [26]),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hF3C0;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[27]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_27))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [27]),
	.datad(\syif.store[27]~input_o ),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hFC30;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\syif.tbCTRL~input_o  & (\syif.store[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_28)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[28]~input_o ),
	.datad(\CPU|DP|PR|Wdata_EX [28]),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hF3C0;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N22
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[29]~input_o ))) # (!\syif.tbCTRL~input_o  & (Wdata_EX_29))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PR|Wdata_EX [29]),
	.datad(\syif.store[29]~input_o ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hFC30;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.tbCTRL~input_o  & (\syif.store[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_30)))

	.dataa(\syif.store[30]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [30]),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hBB88;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\syif.tbCTRL~input_o  & (\syif.store[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((Wdata_EX_31)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[31]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|PR|Wdata_EX [31]),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hDD88;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X1_Y36_N9
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X1_Y36_N13
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X1_Y36_N11
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X1_Y36_N5
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N0
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[1] & (!count[0] & (!count[3] & !count[2])))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[2]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N14
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N8
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[1] & (count[0] & count[2]))))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[2]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N12
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h7878;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N10
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[0] $ (count[1])

	.dataa(gnd),
	.datab(count[0]),
	.datac(count[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h3C3C;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y36_N4
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[1]) # ((count[3]) # (count[2]))))

	.dataa(count[1]),
	.datab(count[3]),
	.datac(count[0]),
	.datad(count[2]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N22
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X65_Y37_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y37_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y37_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11 .lut_mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hA50A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'h88DD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hF3C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hBF80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h0700;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hAAC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hBA10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .lut_mask = 16'h0030;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .lut_mask = 16'hBB42;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .lut_mask = 16'hF0CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hC001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0002;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h2E10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h3CF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .lut_mask = 16'hECA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0008;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~7_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h4040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hF404;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h4400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h3FCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h3CF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .lut_mask = 16'h0429;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hCCCD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'hB9E3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h00AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h0302;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h3320;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .lut_mask = 16'hC0D5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hBA30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFF08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'h01AD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'h1170;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N22
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N8
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y31_N8
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N15
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y0_N1
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N1
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N22
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N8
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N22
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N8
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N22
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y0_N22
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N15
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N15
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N15
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N15
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N8
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N1
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N15
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N8
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N1
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N15
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N22
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N22
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y32_N8
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N15
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N15
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y31_N1
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y0_N15
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N15
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y32_N1
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N22
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N22
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N22
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N15
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N22
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N22
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G0
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G3
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N9
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|halt_reg~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y0_N9
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N9
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X45_Y0_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y29_N16
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N16
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y73_N23
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N2
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N9
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N9
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y30_N9
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y0_N16
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N2
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N23
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N2
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N23
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N23
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N2
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X45_Y0_N16
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N9
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y0_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N23
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y0_N23
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N2
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y31_N16
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h3373;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFB;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hF0AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hA080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N22
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hD2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h0080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h7430;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h22F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hFA0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hA808;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h3300;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFCFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h22AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFEF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hADA8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hA8B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hB9A8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h1C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X10_Y45_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	Result_EX_1,
	pc_1,
	Memwrite_EX,
	MemToReg_EX,
	Result_EX_0,
	pc_0,
	Result_EX_3,
	pc_3,
	Result_EX_2,
	pc_2,
	Result_EX_5,
	pc_5,
	Result_EX_4,
	pc_4,
	Result_EX_7,
	pc_7,
	Result_EX_6,
	pc_6,
	Result_EX_9,
	pc_9,
	Result_EX_8,
	pc_8,
	Result_EX_11,
	pc_11,
	Result_EX_10,
	pc_10,
	Result_EX_13,
	pc_13,
	Result_EX_12,
	pc_12,
	Result_EX_15,
	pc_15,
	Result_EX_14,
	pc_14,
	Result_EX_17,
	pc_17,
	Result_EX_16,
	pc_16,
	Result_EX_19,
	pc_19,
	Result_EX_18,
	pc_18,
	Result_EX_21,
	pc_21,
	Result_EX_20,
	pc_20,
	Result_EX_23,
	pc_23,
	Result_EX_22,
	pc_22,
	Result_EX_25,
	pc_25,
	Result_EX_24,
	pc_24,
	Result_EX_27,
	pc_27,
	Result_EX_26,
	pc_26,
	Result_EX_29,
	pc_29,
	Result_EX_28,
	pc_28,
	Result_EX_31,
	pc_31,
	Result_EX_30,
	pc_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	Wdata_EX_0,
	Wdata_EX_1,
	Wdata_EX_2,
	Wdata_EX_3,
	Wdata_EX_4,
	Wdata_EX_5,
	Wdata_EX_6,
	Wdata_EX_7,
	Wdata_EX_8,
	Wdata_EX_9,
	Wdata_EX_10,
	Wdata_EX_11,
	Wdata_EX_12,
	Wdata_EX_13,
	Wdata_EX_14,
	Wdata_EX_15,
	Wdata_EX_16,
	Wdata_EX_17,
	Wdata_EX_18,
	Wdata_EX_19,
	Wdata_EX_20,
	Wdata_EX_21,
	Wdata_EX_22,
	Wdata_EX_23,
	Wdata_EX_24,
	Wdata_EX_25,
	Wdata_EX_26,
	Wdata_EX_27,
	Wdata_EX_28,
	Wdata_EX_29,
	Wdata_EX_30,
	Wdata_EX_31,
	CLK,
	nRST,
	halt_reg,
	devpor,
	devclrn,
	devoe);
output 	Result_EX_1;
output 	pc_1;
output 	Memwrite_EX;
output 	MemToReg_EX;
output 	Result_EX_0;
output 	pc_0;
output 	Result_EX_3;
output 	pc_3;
output 	Result_EX_2;
output 	pc_2;
output 	Result_EX_5;
output 	pc_5;
output 	Result_EX_4;
output 	pc_4;
output 	Result_EX_7;
output 	pc_7;
output 	Result_EX_6;
output 	pc_6;
output 	Result_EX_9;
output 	pc_9;
output 	Result_EX_8;
output 	pc_8;
output 	Result_EX_11;
output 	pc_11;
output 	Result_EX_10;
output 	pc_10;
output 	Result_EX_13;
output 	pc_13;
output 	Result_EX_12;
output 	pc_12;
output 	Result_EX_15;
output 	pc_15;
output 	Result_EX_14;
output 	pc_14;
output 	Result_EX_17;
output 	pc_17;
output 	Result_EX_16;
output 	pc_16;
output 	Result_EX_19;
output 	pc_19;
output 	Result_EX_18;
output 	pc_18;
output 	Result_EX_21;
output 	pc_21;
output 	Result_EX_20;
output 	pc_20;
output 	Result_EX_23;
output 	pc_23;
output 	Result_EX_22;
output 	pc_22;
output 	Result_EX_25;
output 	pc_25;
output 	Result_EX_24;
output 	pc_24;
output 	Result_EX_27;
output 	pc_27;
output 	Result_EX_26;
output 	pc_26;
output 	Result_EX_29;
output 	pc_29;
output 	Result_EX_28;
output 	pc_28;
output 	Result_EX_31;
output 	pc_31;
output 	Result_EX_30;
output 	pc_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	Wdata_EX_0;
output 	Wdata_EX_1;
output 	Wdata_EX_2;
output 	Wdata_EX_3;
output 	Wdata_EX_4;
output 	Wdata_EX_5;
output 	Wdata_EX_6;
output 	Wdata_EX_7;
output 	Wdata_EX_8;
output 	Wdata_EX_9;
output 	Wdata_EX_10;
output 	Wdata_EX_11;
output 	Wdata_EX_12;
output 	Wdata_EX_13;
output 	Wdata_EX_14;
output 	Wdata_EX_15;
output 	Wdata_EX_16;
output 	Wdata_EX_17;
output 	Wdata_EX_18;
output 	Wdata_EX_19;
output 	Wdata_EX_20;
output 	Wdata_EX_21;
output 	Wdata_EX_22;
output 	Wdata_EX_23;
output 	Wdata_EX_24;
output 	Wdata_EX_25;
output 	Wdata_EX_26;
output 	Wdata_EX_27;
output 	Wdata_EX_28;
output 	Wdata_EX_29;
output 	Wdata_EX_30;
output 	Wdata_EX_31;
input 	CLK;
input 	nRST;
output 	halt_reg;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|always0~0_combout ;


memory_control CC(
	.Memwrite_EX(Memwrite_EX),
	.MemToReg_EX(MemToReg_EX),
	.always0(\CC|always0~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.Result_EX_1(Result_EX_1),
	.pc_1(pc_1),
	.Memwrite_EX(Memwrite_EX),
	.MemToReg_EX(MemToReg_EX),
	.Result_EX_0(Result_EX_0),
	.pc_0(pc_0),
	.Result_EX_3(Result_EX_3),
	.pc_3(pc_3),
	.Result_EX_2(Result_EX_2),
	.pc_2(pc_2),
	.Result_EX_5(Result_EX_5),
	.pc_5(pc_5),
	.Result_EX_4(Result_EX_4),
	.pc_4(pc_4),
	.Result_EX_7(Result_EX_7),
	.pc_7(pc_7),
	.Result_EX_6(Result_EX_6),
	.pc_6(pc_6),
	.Result_EX_9(Result_EX_9),
	.pc_9(pc_9),
	.Result_EX_8(Result_EX_8),
	.pc_8(pc_8),
	.Result_EX_11(Result_EX_11),
	.pc_11(pc_11),
	.Result_EX_10(Result_EX_10),
	.pc_10(pc_10),
	.Result_EX_13(Result_EX_13),
	.pc_13(pc_13),
	.Result_EX_12(Result_EX_12),
	.pc_12(pc_12),
	.Result_EX_15(Result_EX_15),
	.pc_15(pc_15),
	.Result_EX_14(Result_EX_14),
	.pc_14(pc_14),
	.Result_EX_17(Result_EX_17),
	.pc_17(pc_17),
	.Result_EX_16(Result_EX_16),
	.pc_16(pc_16),
	.Result_EX_19(Result_EX_19),
	.pc_19(pc_19),
	.Result_EX_18(Result_EX_18),
	.pc_18(pc_18),
	.Result_EX_21(Result_EX_21),
	.pc_21(pc_21),
	.Result_EX_20(Result_EX_20),
	.pc_20(pc_20),
	.Result_EX_23(Result_EX_23),
	.pc_23(pc_23),
	.Result_EX_22(Result_EX_22),
	.pc_22(pc_22),
	.Result_EX_25(Result_EX_25),
	.pc_25(pc_25),
	.Result_EX_24(Result_EX_24),
	.pc_24(pc_24),
	.Result_EX_27(Result_EX_27),
	.pc_27(pc_27),
	.Result_EX_26(Result_EX_26),
	.pc_26(pc_26),
	.Result_EX_29(Result_EX_29),
	.pc_29(pc_29),
	.Result_EX_28(Result_EX_28),
	.pc_28(pc_28),
	.Result_EX_31(Result_EX_31),
	.pc_31(pc_31),
	.Result_EX_30(Result_EX_30),
	.pc_30(pc_30),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.Wdata_EX_0(Wdata_EX_0),
	.always0(\CC|always0~0_combout ),
	.Wdata_EX_1(Wdata_EX_1),
	.Wdata_EX_2(Wdata_EX_2),
	.Wdata_EX_3(Wdata_EX_3),
	.Wdata_EX_4(Wdata_EX_4),
	.Wdata_EX_5(Wdata_EX_5),
	.Wdata_EX_6(Wdata_EX_6),
	.Wdata_EX_7(Wdata_EX_7),
	.Wdata_EX_8(Wdata_EX_8),
	.Wdata_EX_9(Wdata_EX_9),
	.Wdata_EX_10(Wdata_EX_10),
	.Wdata_EX_11(Wdata_EX_11),
	.Wdata_EX_12(Wdata_EX_12),
	.Wdata_EX_13(Wdata_EX_13),
	.Wdata_EX_14(Wdata_EX_14),
	.Wdata_EX_15(Wdata_EX_15),
	.Wdata_EX_16(Wdata_EX_16),
	.Wdata_EX_17(Wdata_EX_17),
	.Wdata_EX_18(Wdata_EX_18),
	.Wdata_EX_19(Wdata_EX_19),
	.Wdata_EX_20(Wdata_EX_20),
	.Wdata_EX_21(Wdata_EX_21),
	.Wdata_EX_22(Wdata_EX_22),
	.Wdata_EX_23(Wdata_EX_23),
	.Wdata_EX_24(Wdata_EX_24),
	.Wdata_EX_25(Wdata_EX_25),
	.Wdata_EX_26(Wdata_EX_26),
	.Wdata_EX_27(Wdata_EX_27),
	.Wdata_EX_28(Wdata_EX_28),
	.Wdata_EX_29(Wdata_EX_29),
	.Wdata_EX_30(Wdata_EX_30),
	.Wdata_EX_31(Wdata_EX_31),
	.CLK(CLK),
	.nRST(nRST),
	.halt_reg1(halt_reg),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module datapath (
	Result_EX_1,
	pc_1,
	Memwrite_EX,
	MemToReg_EX,
	Result_EX_0,
	pc_0,
	Result_EX_3,
	pc_3,
	Result_EX_2,
	pc_2,
	Result_EX_5,
	pc_5,
	Result_EX_4,
	pc_4,
	Result_EX_7,
	pc_7,
	Result_EX_6,
	pc_6,
	Result_EX_9,
	pc_9,
	Result_EX_8,
	pc_8,
	Result_EX_11,
	pc_11,
	Result_EX_10,
	pc_10,
	Result_EX_13,
	pc_13,
	Result_EX_12,
	pc_12,
	Result_EX_15,
	pc_15,
	Result_EX_14,
	pc_14,
	Result_EX_17,
	pc_17,
	Result_EX_16,
	pc_16,
	Result_EX_19,
	pc_19,
	Result_EX_18,
	pc_18,
	Result_EX_21,
	pc_21,
	Result_EX_20,
	pc_20,
	Result_EX_23,
	pc_23,
	Result_EX_22,
	pc_22,
	Result_EX_25,
	pc_25,
	Result_EX_24,
	pc_24,
	Result_EX_27,
	pc_27,
	Result_EX_26,
	pc_26,
	Result_EX_29,
	pc_29,
	Result_EX_28,
	pc_28,
	Result_EX_31,
	pc_31,
	Result_EX_30,
	pc_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	Wdata_EX_0,
	always0,
	Wdata_EX_1,
	Wdata_EX_2,
	Wdata_EX_3,
	Wdata_EX_4,
	Wdata_EX_5,
	Wdata_EX_6,
	Wdata_EX_7,
	Wdata_EX_8,
	Wdata_EX_9,
	Wdata_EX_10,
	Wdata_EX_11,
	Wdata_EX_12,
	Wdata_EX_13,
	Wdata_EX_14,
	Wdata_EX_15,
	Wdata_EX_16,
	Wdata_EX_17,
	Wdata_EX_18,
	Wdata_EX_19,
	Wdata_EX_20,
	Wdata_EX_21,
	Wdata_EX_22,
	Wdata_EX_23,
	Wdata_EX_24,
	Wdata_EX_25,
	Wdata_EX_26,
	Wdata_EX_27,
	Wdata_EX_28,
	Wdata_EX_29,
	Wdata_EX_30,
	Wdata_EX_31,
	CLK,
	nRST,
	halt_reg1,
	devpor,
	devclrn,
	devoe);
output 	Result_EX_1;
output 	pc_1;
output 	Memwrite_EX;
output 	MemToReg_EX;
output 	Result_EX_0;
output 	pc_0;
output 	Result_EX_3;
output 	pc_3;
output 	Result_EX_2;
output 	pc_2;
output 	Result_EX_5;
output 	pc_5;
output 	Result_EX_4;
output 	pc_4;
output 	Result_EX_7;
output 	pc_7;
output 	Result_EX_6;
output 	pc_6;
output 	Result_EX_9;
output 	pc_9;
output 	Result_EX_8;
output 	pc_8;
output 	Result_EX_11;
output 	pc_11;
output 	Result_EX_10;
output 	pc_10;
output 	Result_EX_13;
output 	pc_13;
output 	Result_EX_12;
output 	pc_12;
output 	Result_EX_15;
output 	pc_15;
output 	Result_EX_14;
output 	pc_14;
output 	Result_EX_17;
output 	pc_17;
output 	Result_EX_16;
output 	pc_16;
output 	Result_EX_19;
output 	pc_19;
output 	Result_EX_18;
output 	pc_18;
output 	Result_EX_21;
output 	pc_21;
output 	Result_EX_20;
output 	pc_20;
output 	Result_EX_23;
output 	pc_23;
output 	Result_EX_22;
output 	pc_22;
output 	Result_EX_25;
output 	pc_25;
output 	Result_EX_24;
output 	pc_24;
output 	Result_EX_27;
output 	pc_27;
output 	Result_EX_26;
output 	pc_26;
output 	Result_EX_29;
output 	pc_29;
output 	Result_EX_28;
output 	pc_28;
output 	Result_EX_31;
output 	pc_31;
output 	Result_EX_30;
output 	pc_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	Wdata_EX_0;
input 	always0;
output 	Wdata_EX_1;
output 	Wdata_EX_2;
output 	Wdata_EX_3;
output 	Wdata_EX_4;
output 	Wdata_EX_5;
output 	Wdata_EX_6;
output 	Wdata_EX_7;
output 	Wdata_EX_8;
output 	Wdata_EX_9;
output 	Wdata_EX_10;
output 	Wdata_EX_11;
output 	Wdata_EX_12;
output 	Wdata_EX_13;
output 	Wdata_EX_14;
output 	Wdata_EX_15;
output 	Wdata_EX_16;
output 	Wdata_EX_17;
output 	Wdata_EX_18;
output 	Wdata_EX_19;
output 	Wdata_EX_20;
output 	Wdata_EX_21;
output 	Wdata_EX_22;
output 	Wdata_EX_23;
output 	Wdata_EX_24;
output 	Wdata_EX_25;
output 	Wdata_EX_26;
output 	Wdata_EX_27;
output 	Wdata_EX_28;
output 	Wdata_EX_29;
output 	Wdata_EX_30;
output 	Wdata_EX_31;
input 	CLK;
input 	nRST;
output 	halt_reg1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \ALU|Add1~62_combout ;
wire \ALU|Add0~42_combout ;
wire \ALU|Add0~44_combout ;
wire \ALU|Add0~46_combout ;
wire \ALU|Add0~48_combout ;
wire \ALU|Add0~50_combout ;
wire \ALU|Add0~52_combout ;
wire \ALU|Add0~54_combout ;
wire \ALU|Add0~56_combout ;
wire \ALU|Add0~58_combout ;
wire \ALU|Add0~60_combout ;
wire \ALU|Add0~62_combout ;
wire \pc_next_branch[2]~0_combout ;
wire \pc_next_branch[8]~12_combout ;
wire \pc_next_branch[16]~28_combout ;
wire \pc_next_branch[17]~30_combout ;
wire \pc_next_branch[18]~32_combout ;
wire \pc_next_branch[20]~36_combout ;
wire \pc_next_branch[29]~55 ;
wire \pc_next_branch[30]~57 ;
wire \pc_next_branch[30]~56_combout ;
wire \pc_next_branch[31]~58_combout ;
wire \PR|halt_MEM~q ;
wire \PR|care_ID~q ;
wire \PR|RegWen_EX~q ;
wire \PR|hazard_Reg_ID~q ;
wire \HZ|always0~0_combout ;
wire \HZ|Equal4~2_combout ;
wire \HZ|Equal4~3_combout ;
wire \PR|Memwrite_ID~q ;
wire \HZ|Equal4~4_combout ;
wire \input_b~0_combout ;
wire \input_b~1_combout ;
wire \PR|MemToReg_MEM~q ;
wire \input_a~56_combout ;
wire \HZ|always0~1_combout ;
wire \PR|RegWen_MEM~q ;
wire \output_RegWen_MEM~0_combout ;
wire \output_RegWen_MEM~1_combout ;
wire \HZ|src2_hazard_t~2_combout ;
wire \input_b~2_combout ;
wire \input_b~3_combout ;
wire \input_b~4_combout ;
wire \input_b~5_combout ;
wire \HZ|always0~2_combout ;
wire \HZ|Equal0~2_combout ;
wire \HZ|Equal0~3_combout ;
wire \input_a~57_combout ;
wire \input_a~58_combout ;
wire \HZ|always0~8_combout ;
wire \HZ|src1_hazard_t~1_combout ;
wire \input_a~59_combout ;
wire \input_a~60_combout ;
wire \input_a~61_combout ;
wire \ALU|out~0_combout ;
wire \input_b~6_combout ;
wire \input_a~62_combout ;
wire \input_b~7_combout ;
wire \input_a~63_combout ;
wire \input_b~8_combout ;
wire \input_b~9_combout ;
wire \input_a~64_combout ;
wire \input_b~10_combout ;
wire \input_a~65_combout ;
wire \input_b~11_combout ;
wire \input_b~12_combout ;
wire \input_a~66_combout ;
wire \input_b~13_combout ;
wire \input_a~67_combout ;
wire \input_b~14_combout ;
wire \input_b~15_combout ;
wire \input_a~68_combout ;
wire \input_b~16_combout ;
wire \input_a~69_combout ;
wire \input_b~17_combout ;
wire \input_b~18_combout ;
wire \input_a~70_combout ;
wire \input_b~19_combout ;
wire \input_a~71_combout ;
wire \input_b~20_combout ;
wire \input_b~21_combout ;
wire \input_a~72_combout ;
wire \input_b~22_combout ;
wire \input_a~73_combout ;
wire \input_b~23_combout ;
wire \input_b~24_combout ;
wire \input_a~74_combout ;
wire \input_b~25_combout ;
wire \input_a~75_combout ;
wire \input_b~26_combout ;
wire \input_b~27_combout ;
wire \input_a~76_combout ;
wire \input_b~28_combout ;
wire \input_a~77_combout ;
wire \input_b~29_combout ;
wire \input_b~30_combout ;
wire \input_a~78_combout ;
wire \input_b~31_combout ;
wire \input_a~79_combout ;
wire \input_b~32_combout ;
wire \input_b~33_combout ;
wire \input_a~80_combout ;
wire \input_b~34_combout ;
wire \input_a~81_combout ;
wire \input_b~35_combout ;
wire \input_b~36_combout ;
wire \input_a~82_combout ;
wire \input_b~37_combout ;
wire \input_a~83_combout ;
wire \input_b~38_combout ;
wire \input_b~39_combout ;
wire \input_a~84_combout ;
wire \input_b~40_combout ;
wire \input_a~85_combout ;
wire \input_b~41_combout ;
wire \input_b~42_combout ;
wire \input_a~86_combout ;
wire \input_b~43_combout ;
wire \input_a~87_combout ;
wire \input_b~44_combout ;
wire \input_b~45_combout ;
wire \input_a~88_combout ;
wire \input_b~46_combout ;
wire \input_a~89_combout ;
wire \input_b~47_combout ;
wire \input_b~48_combout ;
wire \input_a~90_combout ;
wire \input_b~49_combout ;
wire \input_a~91_combout ;
wire \input_b~50_combout ;
wire \input_b~51_combout ;
wire \input_a~92_combout ;
wire \input_b~52_combout ;
wire \input_a~93_combout ;
wire \input_b~53_combout ;
wire \input_b~54_combout ;
wire \input_a~94_combout ;
wire \input_b~55_combout ;
wire \input_a~95_combout ;
wire \input_b~56_combout ;
wire \input_b~57_combout ;
wire \input_a~96_combout ;
wire \input_b~58_combout ;
wire \input_b~59_combout ;
wire \input_a~97_combout ;
wire \input_a~98_combout ;
wire \input_a~99_combout ;
wire \input_b~60_combout ;
wire \input_b~61_combout ;
wire \input_a~100_combout ;
wire \input_a~101_combout ;
wire \input_a~102_combout ;
wire \input_b~62_combout ;
wire \input_b~63_combout ;
wire \input_a~103_combout ;
wire \input_a~104_combout ;
wire \input_a~105_combout ;
wire \input_b~64_combout ;
wire \input_b~65_combout ;
wire \input_a~106_combout ;
wire \input_a~107_combout ;
wire \input_a~108_combout ;
wire \input_b~66_combout ;
wire \input_b~67_combout ;
wire \input_a~109_combout ;
wire \input_a~110_combout ;
wire \input_a~111_combout ;
wire \input_b~68_combout ;
wire \input_b~69_combout ;
wire \input_a~112_combout ;
wire \input_a~113_combout ;
wire \input_a~114_combout ;
wire \input_b~70_combout ;
wire \input_b~71_combout ;
wire \input_a~115_combout ;
wire \input_a~116_combout ;
wire \input_a~117_combout ;
wire \input_b~72_combout ;
wire \input_b~73_combout ;
wire \input_a~118_combout ;
wire \input_a~119_combout ;
wire \input_a~120_combout ;
wire \input_b~74_combout ;
wire \input_b~75_combout ;
wire \input_a~121_combout ;
wire \input_a~122_combout ;
wire \input_a~123_combout ;
wire \input_b~76_combout ;
wire \input_b~77_combout ;
wire \input_a~124_combout ;
wire \input_a~125_combout ;
wire \input_a~126_combout ;
wire \input_b~78_combout ;
wire \input_b~79_combout ;
wire \input_a~127_combout ;
wire \input_a~128_combout ;
wire \input_a~129_combout ;
wire \input_b~80_combout ;
wire \input_b~81_combout ;
wire \input_a~130_combout ;
wire \input_a~131_combout ;
wire \input_b~82_combout ;
wire \input_b~83_combout ;
wire \input_a~133_combout ;
wire \input_a~134_combout ;
wire \input_b~84_combout ;
wire \input_b~85_combout ;
wire \input_a~136_combout ;
wire \input_a~137_combout ;
wire \ALU|Equal0~0_combout ;
wire \ALU|Equal0~5_combout ;
wire \ALU|Equal0~6_combout ;
wire \HZ|src2_hazard_t~3_combout ;
wire \ALU|Selector30~7_combout ;
wire \halt_reg~10_combout ;
wire \ALU|Selector28~10_combout ;
wire \ALU|Selector3~11_combout ;
wire \ALU|Selector22~9_combout ;
wire \ALU|Selector2~8_combout ;
wire \ALU|Selector27~8_combout ;
wire \ALU|Selector25~7_combout ;
wire \input_b~86_combout ;
wire \ALU|Selector24~8_combout ;
wire \ALU|Selector26~7_combout ;
wire \ALU|Selector4~7_combout ;
wire \ALU|Selector16~10_combout ;
wire \ALU|Selector7~12_combout ;
wire \ALU|Selector6~6_combout ;
wire \ALU|Selector29~10_combout ;
wire \ALU|Selector15~14_combout ;
wire \ALU|Selector5~6_combout ;
wire \ALU|Selector31~11_combout ;
wire \ALU|Selector11~9_combout ;
wire \ALU|Selector10~8_combout ;
wire \ALU|Selector21~9_combout ;
wire \ALU|Selector20~8_combout ;
wire \ALU|Selector9~8_combout ;
wire \ALU|Selector8~8_combout ;
wire \ALU|Selector14~7_combout ;
wire \ALU|Selector13~7_combout ;
wire \ALU|Selector12~7_combout ;
wire \ALU|Selector23~10_combout ;
wire \ALU|Selector19~9_combout ;
wire \ALU|Selector18~8_combout ;
wire \ALU|Selector17~7_combout ;
wire \ALU|Selector0~28_combout ;
wire \ALU|Selector1~11_combout ;
wire \ALU|Equal11~11_combout ;
wire \input_a~138_combout ;
wire \pc_next[3]~6_combout ;
wire \input_a~139_combout ;
wire \pc_next[5]~15_combout ;
wire \pc_next[7]~23_combout ;
wire \pc_next[6]~27_combout ;
wire \pc_next[19]~71_combout ;
wire \pc_next[19]~72_combout ;
wire \pc_next[21]~79_combout ;
wire \pc_next[21]~80_combout ;
wire \pc_next[27]~103_combout ;
wire \pc[29]~29_combout ;
wire \pc_next[28]~114_combout ;
wire \CU|Selector14~0_combout ;
wire \HZ|src2_hazard_t~4_combout ;
wire \CU|Selector11~0_combout ;
wire \CU|WideOr4~0_combout ;
wire \CU|WideOr4~1_combout ;
wire \CU|input_hazard_Reg_ID~0_combout ;
wire \CU|WideOr21~0_combout ;
wire \Equal20~0_combout ;
wire \CU|Selector14~2_combout ;
wire \CU|WideOr21~2_combout ;
wire \CU|WideOr21~3_combout ;
wire \RF|rfif.rdat2[31]~20_combout ;
wire \CU|WideOr14~0_combout ;
wire \RF|rfif.rdat1[31]~9_combout ;
wire \RF|rfif.rdat1[31]~19_combout ;
wire \RF|WideOr0~0_combout ;
wire \CU|WideOr6~0_combout ;
wire \CU|WideOr6~1_combout ;
wire \RF|rfif.rdat1[30]~29_combout ;
wire \RF|rfif.rdat1[30]~39_combout ;
wire \RF|rfif.rdat2[30]~41_combout ;
wire \RF|rfif.rdat1[29]~49_combout ;
wire \RF|rfif.rdat1[29]~59_combout ;
wire \RF|rfif.rdat2[29]~62_combout ;
wire \RF|rfif.rdat1[28]~69_combout ;
wire \RF|rfif.rdat1[28]~79_combout ;
wire \RF|rfif.rdat2[28]~83_combout ;
wire \RF|rfif.rdat1[27]~89_combout ;
wire \RF|rfif.rdat1[27]~99_combout ;
wire \RF|rfif.rdat2[27]~104_combout ;
wire \RF|rfif.rdat1[26]~109_combout ;
wire \RF|rfif.rdat1[26]~119_combout ;
wire \RF|rfif.rdat2[26]~125_combout ;
wire \RF|rfif.rdat1[25]~129_combout ;
wire \RF|rfif.rdat1[25]~139_combout ;
wire \RF|rfif.rdat2[25]~146_combout ;
wire \RF|rfif.rdat1[24]~149_combout ;
wire \RF|rfif.rdat1[24]~159_combout ;
wire \RF|rfif.rdat2[24]~167_combout ;
wire \RF|rfif.rdat1[23]~169_combout ;
wire \RF|rfif.rdat1[23]~179_combout ;
wire \RF|rfif.rdat2[23]~188_combout ;
wire \RF|rfif.rdat1[22]~189_combout ;
wire \RF|rfif.rdat1[22]~199_combout ;
wire \RF|rfif.rdat2[22]~209_combout ;
wire \RF|rfif.rdat1[21]~209_combout ;
wire \RF|rfif.rdat1[21]~219_combout ;
wire \RF|rfif.rdat2[21]~230_combout ;
wire \RF|rfif.rdat1[20]~229_combout ;
wire \RF|rfif.rdat1[20]~239_combout ;
wire \RF|rfif.rdat2[20]~251_combout ;
wire \RF|rfif.rdat1[19]~249_combout ;
wire \RF|rfif.rdat1[19]~259_combout ;
wire \RF|rfif.rdat2[19]~272_combout ;
wire \RF|rfif.rdat1[18]~269_combout ;
wire \RF|rfif.rdat1[18]~279_combout ;
wire \RF|rfif.rdat2[18]~293_combout ;
wire \RF|rfif.rdat1[17]~289_combout ;
wire \RF|rfif.rdat1[17]~299_combout ;
wire \RF|rfif.rdat2[17]~314_combout ;
wire \RF|rfif.rdat1[16]~309_combout ;
wire \RF|rfif.rdat1[16]~319_combout ;
wire \RF|rfif.rdat2[16]~335_combout ;
wire \RF|rfif.rdat1[15]~329_combout ;
wire \RF|rfif.rdat1[15]~339_combout ;
wire \Equal0~0_combout ;
wire \RF|rfif.rdat2[15]~356_combout ;
wire \RF|rfif.rdat1[14]~349_combout ;
wire \RF|rfif.rdat1[14]~359_combout ;
wire \RF|rfif.rdat2[14]~377_combout ;
wire \RF|rfif.rdat2[13]~398_combout ;
wire \RF|rfif.rdat1[13]~369_combout ;
wire \RF|rfif.rdat1[13]~379_combout ;
wire \RF|rfif.rdat2[12]~419_combout ;
wire \RF|rfif.rdat1[12]~389_combout ;
wire \RF|rfif.rdat1[12]~399_combout ;
wire \RF|rfif.rdat2[11]~440_combout ;
wire \RF|rfif.rdat1[11]~409_combout ;
wire \RF|rfif.rdat1[11]~419_combout ;
wire \RF|rfif.rdat2[10]~461_combout ;
wire \RF|rfif.rdat1[10]~429_combout ;
wire \RF|rfif.rdat1[10]~439_combout ;
wire \RF|rfif.rdat2[9]~482_combout ;
wire \RF|rfif.rdat1[9]~449_combout ;
wire \RF|rfif.rdat1[9]~459_combout ;
wire \RF|rfif.rdat2[8]~503_combout ;
wire \RF|rfif.rdat1[8]~469_combout ;
wire \RF|rfif.rdat1[8]~479_combout ;
wire \RF|rfif.rdat2[7]~524_combout ;
wire \RF|rfif.rdat1[7]~489_combout ;
wire \RF|rfif.rdat1[7]~499_combout ;
wire \RF|rfif.rdat2[6]~545_combout ;
wire \RF|rfif.rdat1[6]~509_combout ;
wire \RF|rfif.rdat1[6]~519_combout ;
wire \RF|rfif.rdat2[5]~566_combout ;
wire \RF|rfif.rdat1[5]~529_combout ;
wire \RF|rfif.rdat1[5]~539_combout ;
wire \RF|rfif.rdat2[4]~587_combout ;
wire \Equal2~0_combout ;
wire \input_ALUSrc2_ID~0_combout ;
wire \input_ALUSrc2_ID~1_combout ;
wire \input_ALUSrc2_ID~2_combout ;
wire \input_ALUSrc2_ID~3_combout ;
wire \RF|rfif.rdat1[4]~549_combout ;
wire \RF|rfif.rdat1[4]~559_combout ;
wire \RF|rfif.rdat2[3]~608_combout ;
wire \input_ALUSrc2_ID~4_combout ;
wire \input_ALUSrc2_ID~5_combout ;
wire \RF|rfif.rdat1[3]~569_combout ;
wire \RF|rfif.rdat1[3]~579_combout ;
wire \RF|rfif.rdat2[2]~629_combout ;
wire \input_ALUSrc2_ID~6_combout ;
wire \input_ALUSrc2_ID~7_combout ;
wire \RF|rfif.rdat1[2]~589_combout ;
wire \RF|rfif.rdat1[2]~599_combout ;
wire \RF|rfif.rdat2[1]~650_combout ;
wire \input_ALUSrc2_ID~8_combout ;
wire \input_ALUSrc2_ID~9_combout ;
wire \RF|rfif.rdat1[1]~609_combout ;
wire \RF|rfif.rdat1[1]~619_combout ;
wire \RF|rfif.rdat2[0]~671_combout ;
wire \input_ALUSrc2_ID~10_combout ;
wire \input_ALUSrc2_ID~11_combout ;
wire \RF|rfif.rdat1[0]~629_combout ;
wire \RF|rfif.rdat1[0]~639_combout ;
wire \Equal27~0_combout ;
wire \CU|WideOr33~0_combout ;
wire \CU|Decoder0~1_combout ;
wire \CU|WideOr11~0_combout ;
wire \input_a~141_combout ;
wire \input_a~142_combout ;
wire \input_a~143_combout ;
wire \input_a~145_combout ;
wire \input_a~152_combout ;
wire \input_a~155_combout ;
wire \input_a~157_combout ;
wire \input_a~162_combout ;
wire \input_a~163_combout ;
wire \input_a~165_combout ;
wire \input_a~166_combout ;
wire \Equal8~0_combout ;
wire \Equal24~0_combout ;
wire \Equal8~1_combout ;
wire \pc[0]~37_combout ;
wire \pc_next~0_combout ;
wire \input_a~132_combout ;
wire \Equal22~0_combout ;
wire \pc[0]~25_combout ;
wire \pc_next~1_combout ;
wire \pc_next~2_combout ;
wire \branch~0_combout ;
wire \pc[1]~26_combout ;
wire \pc[1]~27_combout ;
wire \pc[0]~24_combout ;
wire \pc[0]~33_combout ;
wire \pc_next~3_combout ;
wire \input_a~135_combout ;
wire \pc_next~4_combout ;
wire \pc_next~5_combout ;
wire \pc_next_plus4[2]~1 ;
wire \pc_next_plus4[3]~2_combout ;
wire \pc_next_branch[2]~1 ;
wire \pc_next_branch[3]~2_combout ;
wire \pc[22]~38_combout ;
wire \pc_next[3]~7_combout ;
wire \pc[22]~28_combout ;
wire \pc_next[3]~8_combout ;
wire \pc_next[27]~9_combout ;
wire \pc_next[3]~10_combout ;
wire \PC_enable~2_combout ;
wire \pc[22]~34_combout ;
wire \pc_next[2]~11_combout ;
wire \pc_next[2]~12_combout ;
wire \pc_next[2]~13_combout ;
wire \pc_next_plus4[2]~0_combout ;
wire \pc_next[2]~14_combout ;
wire \pc_next_plus4[3]~3 ;
wire \pc_next_plus4[4]~5 ;
wire \pc_next_plus4[5]~6_combout ;
wire \pc_next[5]~16_combout ;
wire \pc_next_branch[3]~3 ;
wire \pc_next_branch[4]~5 ;
wire \pc_next_branch[5]~6_combout ;
wire \pc_next[5]~17_combout ;
wire \pc_next[5]~18_combout ;
wire \pc_next_plus4[4]~4_combout ;
wire \input_a~140_combout ;
wire \pc_next[4]~19_combout ;
wire \pc_next[4]~20_combout ;
wire \pc_next_branch[4]~4_combout ;
wire \pc_next[4]~21_combout ;
wire \pc_next[4]~22_combout ;
wire \pc_next_branch[5]~7 ;
wire \pc_next_branch[6]~9 ;
wire \pc_next_branch[7]~10_combout ;
wire \pc_next[7]~24_combout ;
wire \pc_next[7]~25_combout ;
wire \pc_next_plus4[5]~7 ;
wire \pc_next_plus4[6]~9 ;
wire \pc_next_plus4[7]~10_combout ;
wire \pc_next[7]~26_combout ;
wire \pc_next_plus4[6]~8_combout ;
wire \pc_next_branch[6]~8_combout ;
wire \input_a~144_combout ;
wire \pc_next[6]~28_combout ;
wire \pc_next[6]~29_combout ;
wire \pc_next[6]~30_combout ;
wire \pc_next[9]~31_combout ;
wire \pc_next[9]~32_combout ;
wire \pc_next_branch[7]~11 ;
wire \pc_next_branch[8]~13 ;
wire \pc_next_branch[9]~14_combout ;
wire \pc_next[9]~33_combout ;
wire \pc_next_plus4[7]~11 ;
wire \pc_next_plus4[8]~13 ;
wire \pc_next_plus4[9]~14_combout ;
wire \pc_next[9]~34_combout ;
wire \pc_next[8]~35_combout ;
wire \input_a~146_combout ;
wire \pc_next[8]~36_combout ;
wire \pc_next[8]~37_combout ;
wire \pc_next_plus4[8]~12_combout ;
wire \pc_next[8]~38_combout ;
wire \pc_next_plus4[9]~15 ;
wire \pc_next_plus4[10]~17 ;
wire \pc_next_plus4[11]~18_combout ;
wire \input_a~147_combout ;
wire \pc_next[11]~39_combout ;
wire \pc_next[11]~40_combout ;
wire \pc_next_branch[9]~15 ;
wire \pc_next_branch[10]~17 ;
wire \pc_next_branch[11]~18_combout ;
wire \pc_next[11]~41_combout ;
wire \pc_next[11]~42_combout ;
wire \pc_next_plus4[10]~16_combout ;
wire \pc_next_branch[10]~16_combout ;
wire \pc_next[10]~43_combout ;
wire \input_a~148_combout ;
wire \pc_next[10]~44_combout ;
wire \pc_next[10]~45_combout ;
wire \pc_next[10]~46_combout ;
wire \pc_next_plus4[11]~19 ;
wire \pc_next_plus4[12]~21 ;
wire \pc_next_plus4[13]~22_combout ;
wire \pc_next_branch[11]~19 ;
wire \pc_next_branch[12]~21 ;
wire \pc_next_branch[13]~22_combout ;
wire \input_a~149_combout ;
wire \pc_next[13]~47_combout ;
wire \pc_next[13]~48_combout ;
wire \pc_next[13]~49_combout ;
wire \pc_next[13]~50_combout ;
wire \input_a~150_combout ;
wire \pc_next[12]~51_combout ;
wire \pc_next[12]~52_combout ;
wire \pc_next_branch[12]~20_combout ;
wire \pc_next[12]~53_combout ;
wire \pc_next_plus4[12]~20_combout ;
wire \pc_next[12]~54_combout ;
wire \input_a~151_combout ;
wire \pc_next[15]~55_combout ;
wire \pc_next[15]~56_combout ;
wire \pc_next_branch[13]~23 ;
wire \pc_next_branch[14]~25 ;
wire \pc_next_branch[15]~26_combout ;
wire \pc_next[15]~57_combout ;
wire \pc_next_plus4[13]~23 ;
wire \pc_next_plus4[14]~25 ;
wire \pc_next_plus4[15]~26_combout ;
wire \pc_next[15]~58_combout ;
wire \pc_next_plus4[14]~24_combout ;
wire \pc_next[14]~59_combout ;
wire \pc_next[14]~60_combout ;
wire \pc_next_branch[14]~24_combout ;
wire \pc_next[14]~61_combout ;
wire \pc_next[14]~62_combout ;
wire \pc_next_plus4[15]~27 ;
wire \pc_next_plus4[16]~29 ;
wire \pc_next_plus4[17]~30_combout ;
wire \input_a~153_combout ;
wire \pc_next[17]~63_combout ;
wire \pc_next[17]~64_combout ;
wire \pc_next[17]~65_combout ;
wire \pc_next[17]~66_combout ;
wire \pc_next_plus4[16]~28_combout ;
wire \input_a~154_combout ;
wire \pc_next[16]~67_combout ;
wire \pc_next[16]~68_combout ;
wire \pc_next[16]~69_combout ;
wire \pc_next[16]~70_combout ;
wire \pc_next_branch[15]~27 ;
wire \pc_next_branch[16]~29 ;
wire \pc_next_branch[17]~31 ;
wire \pc_next_branch[18]~33 ;
wire \pc_next_branch[19]~34_combout ;
wire \pc_next[19]~73_combout ;
wire \pc_next_plus4[17]~31 ;
wire \pc_next_plus4[18]~33 ;
wire \pc_next_plus4[19]~34_combout ;
wire \pc_next[19]~74_combout ;
wire \pc_next_plus4[18]~32_combout ;
wire \pc_next[18]~75_combout ;
wire \input_a~156_combout ;
wire \pc_next[18]~76_combout ;
wire \pc_next[18]~77_combout ;
wire \pc_next[18]~78_combout ;
wire \pc_next_branch[19]~35 ;
wire \pc_next_branch[20]~37 ;
wire \pc_next_branch[21]~38_combout ;
wire \pc_next[21]~81_combout ;
wire \pc_next_plus4[19]~35 ;
wire \pc_next_plus4[20]~37 ;
wire \pc_next_plus4[21]~38_combout ;
wire \pc_next[21]~82_combout ;
wire \pc_next[20]~83_combout ;
wire \input_a~158_combout ;
wire \pc_next[20]~84_combout ;
wire \pc_next[20]~85_combout ;
wire \pc_next_plus4[20]~36_combout ;
wire \pc_next[20]~86_combout ;
wire \input_a~159_combout ;
wire \pc_next[23]~87_combout ;
wire \pc_next[23]~88_combout ;
wire \pc_next_branch[21]~39 ;
wire \pc_next_branch[22]~41 ;
wire \pc_next_branch[23]~42_combout ;
wire \pc_next[23]~89_combout ;
wire \pc_next_plus4[21]~39 ;
wire \pc_next_plus4[22]~41 ;
wire \pc_next_plus4[23]~42_combout ;
wire \pc_next[23]~90_combout ;
wire \pc_next_branch[22]~40_combout ;
wire \input_a~160_combout ;
wire \pc_next[22]~91_combout ;
wire \pc_next[22]~92_combout ;
wire \pc_next[22]~93_combout ;
wire \pc_next_plus4[22]~40_combout ;
wire \pc_next[22]~94_combout ;
wire \input_a~161_combout ;
wire \pc_next[25]~95_combout ;
wire \pc_next[25]~96_combout ;
wire \pc_next_branch[23]~43 ;
wire \pc_next_branch[24]~45 ;
wire \pc_next_branch[25]~46_combout ;
wire \pc_next[25]~97_combout ;
wire \pc_next_plus4[23]~43 ;
wire \pc_next_plus4[24]~45 ;
wire \pc_next_plus4[25]~46_combout ;
wire \pc_next[25]~98_combout ;
wire \pc_next[24]~99_combout ;
wire \pc_next[24]~100_combout ;
wire \pc_next_branch[24]~44_combout ;
wire \pc_next[24]~101_combout ;
wire \pc_next_plus4[24]~44_combout ;
wire \pc_next[24]~102_combout ;
wire \pc_next_plus4[25]~47 ;
wire \pc_next_plus4[26]~49 ;
wire \pc_next_plus4[27]~50_combout ;
wire \pc_next[27]~104_combout ;
wire \pc_next_branch[25]~47 ;
wire \pc_next_branch[26]~49 ;
wire \pc_next_branch[27]~50_combout ;
wire \pc_next[27]~105_combout ;
wire \pc_next[27]~106_combout ;
wire \pc_next_plus4[26]~48_combout ;
wire \pc_next_branch[26]~48_combout ;
wire \input_a~164_combout ;
wire \pc_next[26]~107_combout ;
wire \pc_next[26]~108_combout ;
wire \pc_next[26]~109_combout ;
wire \pc_next[26]~110_combout ;
wire \pc[29]~35_combout ;
wire \Equal23~0_combout ;
wire \pc[29]~31_combout ;
wire \pc[29]~30_combout ;
wire \pc_next[29]~111_combout ;
wire \pc_next_branch[27]~51 ;
wire \pc_next_branch[28]~53 ;
wire \pc_next_branch[29]~54_combout ;
wire \pc_next[29]~112_combout ;
wire \pc_next_plus4[27]~51 ;
wire \pc_next_plus4[28]~53 ;
wire \pc_next_plus4[29]~54_combout ;
wire \pc[29]~36_combout ;
wire \pc_next[29]~113_combout ;
wire \pc[31]~32_combout ;
wire \pc_next_plus4[28]~52_combout ;
wire \pc_next_branch[28]~52_combout ;
wire \pc_next[28]~115_combout ;
wire \pc_next[28]~116_combout ;
wire \input_a~167_combout ;
wire \pc_next[31]~117_combout ;
wire \pc_next[31]~118_combout ;
wire \pc_next_plus4[29]~55 ;
wire \pc_next_plus4[30]~57 ;
wire \pc_next_plus4[31]~58_combout ;
wire \pc_next[31]~119_combout ;
wire \input_a~168_combout ;
wire \pc_next[30]~120_combout ;
wire \pc_next[30]~121_combout ;
wire \pc_next_plus4[30]~56_combout ;
wire \pc_next[30]~122_combout ;
wire \halt_reg~_Duplicate_1_q ;
wire \halt_reg~0_combout ;
wire \halt_reg~1_combout ;
wire \halt_reg~2_combout ;
wire \halt_reg~3_combout ;
wire \halt_reg~4_combout ;
wire \halt_reg~5_combout ;
wire \halt_reg~6_combout ;
wire \halt_reg~7_combout ;
wire \halt_reg~8_combout ;
wire \halt_reg~9_combout ;
wire [31:0] \PR|nextPC_ID ;
wire [2:0] \PR|jump_ID ;
wire [4:0] \PR|RegDst_MEM ;
wire [4:0] \PR|RegDst_EX ;
wire [31:0] \PR|ReadData_MEM ;
wire [31:0] \PR|Instr_IF ;
wire [31:0] \PR|Instr_ID ;
wire [31:0] \PR|CalcData_MEM ;
wire [31:0] \PR|ALUSrc2_ID ;
wire [31:0] \PR|ALUSrc1_ID ;
wire [3:0] \PR|ALUOP_ID ;


register_file RF(
	.input_a(\input_a~56_combout ),
	.RegWen_MEM(\PR|RegWen_MEM~q ),
	.RegDst_MEM_0(\PR|RegDst_MEM [0]),
	.RegDst_MEM_1(\PR|RegDst_MEM [1]),
	.RegDst_MEM_4(\PR|RegDst_MEM [4]),
	.RegDst_MEM_3(\PR|RegDst_MEM [3]),
	.RegDst_MEM_2(\PR|RegDst_MEM [2]),
	.input_b(\input_b~7_combout ),
	.input_b1(\input_b~10_combout ),
	.input_b2(\input_b~13_combout ),
	.input_b3(\input_b~16_combout ),
	.input_b4(\input_b~19_combout ),
	.input_b5(\input_b~22_combout ),
	.input_b6(\input_b~25_combout ),
	.input_b7(\input_b~28_combout ),
	.input_b8(\input_b~31_combout ),
	.input_b9(\input_b~34_combout ),
	.input_b10(\input_b~37_combout ),
	.input_b11(\input_b~40_combout ),
	.input_b12(\input_b~43_combout ),
	.input_b13(\input_b~46_combout ),
	.input_b14(\input_b~49_combout ),
	.input_b15(\input_b~52_combout ),
	.input_b16(\input_b~55_combout ),
	.input_a1(\input_a~96_combout ),
	.input_a2(\input_a~99_combout ),
	.input_a3(\input_a~102_combout ),
	.input_a4(\input_a~105_combout ),
	.input_a5(\input_a~108_combout ),
	.input_a6(\input_a~111_combout ),
	.input_a7(\input_a~114_combout ),
	.input_a8(\input_a~117_combout ),
	.input_a9(\input_a~120_combout ),
	.input_a10(\input_a~123_combout ),
	.input_a11(\input_a~126_combout ),
	.input_a12(\input_a~129_combout ),
	.input_a13(\input_a~132_combout ),
	.input_a14(\input_a~135_combout ),
	.Instr_IF_16(\PR|Instr_IF [16]),
	.Instr_IF_17(\PR|Instr_IF [17]),
	.Instr_IF_18(\PR|Instr_IF [18]),
	.Instr_IF_19(\PR|Instr_IF [19]),
	.Instr_IF_20(\PR|Instr_IF [20]),
	.rfifrdat2_31(\RF|rfif.rdat2[31]~20_combout ),
	.Instr_IF_21(\PR|Instr_IF [21]),
	.Instr_IF_22(\PR|Instr_IF [22]),
	.Instr_IF_24(\PR|Instr_IF [24]),
	.Instr_IF_25(\PR|Instr_IF [25]),
	.Instr_IF_23(\PR|Instr_IF [23]),
	.rfifrdat1_31(\RF|rfif.rdat1[31]~9_combout ),
	.rfifrdat1_311(\RF|rfif.rdat1[31]~19_combout ),
	.WideOr0(\RF|WideOr0~0_combout ),
	.rfifrdat1_30(\RF|rfif.rdat1[30]~29_combout ),
	.rfifrdat1_301(\RF|rfif.rdat1[30]~39_combout ),
	.rfifrdat2_30(\RF|rfif.rdat2[30]~41_combout ),
	.rfifrdat1_29(\RF|rfif.rdat1[29]~49_combout ),
	.rfifrdat1_291(\RF|rfif.rdat1[29]~59_combout ),
	.rfifrdat2_29(\RF|rfif.rdat2[29]~62_combout ),
	.rfifrdat1_28(\RF|rfif.rdat1[28]~69_combout ),
	.rfifrdat1_281(\RF|rfif.rdat1[28]~79_combout ),
	.rfifrdat2_28(\RF|rfif.rdat2[28]~83_combout ),
	.rfifrdat1_27(\RF|rfif.rdat1[27]~89_combout ),
	.rfifrdat1_271(\RF|rfif.rdat1[27]~99_combout ),
	.rfifrdat2_27(\RF|rfif.rdat2[27]~104_combout ),
	.rfifrdat1_26(\RF|rfif.rdat1[26]~109_combout ),
	.rfifrdat1_261(\RF|rfif.rdat1[26]~119_combout ),
	.rfifrdat2_26(\RF|rfif.rdat2[26]~125_combout ),
	.rfifrdat1_25(\RF|rfif.rdat1[25]~129_combout ),
	.rfifrdat1_251(\RF|rfif.rdat1[25]~139_combout ),
	.rfifrdat2_25(\RF|rfif.rdat2[25]~146_combout ),
	.rfifrdat1_24(\RF|rfif.rdat1[24]~149_combout ),
	.rfifrdat1_241(\RF|rfif.rdat1[24]~159_combout ),
	.rfifrdat2_24(\RF|rfif.rdat2[24]~167_combout ),
	.rfifrdat1_23(\RF|rfif.rdat1[23]~169_combout ),
	.rfifrdat1_231(\RF|rfif.rdat1[23]~179_combout ),
	.rfifrdat2_23(\RF|rfif.rdat2[23]~188_combout ),
	.rfifrdat1_22(\RF|rfif.rdat1[22]~189_combout ),
	.rfifrdat1_221(\RF|rfif.rdat1[22]~199_combout ),
	.rfifrdat2_22(\RF|rfif.rdat2[22]~209_combout ),
	.rfifrdat1_21(\RF|rfif.rdat1[21]~209_combout ),
	.rfifrdat1_211(\RF|rfif.rdat1[21]~219_combout ),
	.rfifrdat2_21(\RF|rfif.rdat2[21]~230_combout ),
	.rfifrdat1_20(\RF|rfif.rdat1[20]~229_combout ),
	.rfifrdat1_201(\RF|rfif.rdat1[20]~239_combout ),
	.rfifrdat2_20(\RF|rfif.rdat2[20]~251_combout ),
	.rfifrdat1_19(\RF|rfif.rdat1[19]~249_combout ),
	.rfifrdat1_191(\RF|rfif.rdat1[19]~259_combout ),
	.rfifrdat2_19(\RF|rfif.rdat2[19]~272_combout ),
	.rfifrdat1_18(\RF|rfif.rdat1[18]~269_combout ),
	.rfifrdat1_181(\RF|rfif.rdat1[18]~279_combout ),
	.rfifrdat2_18(\RF|rfif.rdat2[18]~293_combout ),
	.rfifrdat1_17(\RF|rfif.rdat1[17]~289_combout ),
	.rfifrdat1_171(\RF|rfif.rdat1[17]~299_combout ),
	.rfifrdat2_17(\RF|rfif.rdat2[17]~314_combout ),
	.rfifrdat1_16(\RF|rfif.rdat1[16]~309_combout ),
	.rfifrdat1_161(\RF|rfif.rdat1[16]~319_combout ),
	.rfifrdat2_16(\RF|rfif.rdat2[16]~335_combout ),
	.rfifrdat1_15(\RF|rfif.rdat1[15]~329_combout ),
	.rfifrdat1_151(\RF|rfif.rdat1[15]~339_combout ),
	.rfifrdat2_15(\RF|rfif.rdat2[15]~356_combout ),
	.rfifrdat1_14(\RF|rfif.rdat1[14]~349_combout ),
	.rfifrdat1_141(\RF|rfif.rdat1[14]~359_combout ),
	.rfifrdat2_14(\RF|rfif.rdat2[14]~377_combout ),
	.rfifrdat2_13(\RF|rfif.rdat2[13]~398_combout ),
	.rfifrdat1_13(\RF|rfif.rdat1[13]~369_combout ),
	.rfifrdat1_131(\RF|rfif.rdat1[13]~379_combout ),
	.rfifrdat2_12(\RF|rfif.rdat2[12]~419_combout ),
	.rfifrdat1_12(\RF|rfif.rdat1[12]~389_combout ),
	.rfifrdat1_121(\RF|rfif.rdat1[12]~399_combout ),
	.rfifrdat2_11(\RF|rfif.rdat2[11]~440_combout ),
	.rfifrdat1_11(\RF|rfif.rdat1[11]~409_combout ),
	.rfifrdat1_111(\RF|rfif.rdat1[11]~419_combout ),
	.rfifrdat2_10(\RF|rfif.rdat2[10]~461_combout ),
	.rfifrdat1_10(\RF|rfif.rdat1[10]~429_combout ),
	.rfifrdat1_101(\RF|rfif.rdat1[10]~439_combout ),
	.rfifrdat2_9(\RF|rfif.rdat2[9]~482_combout ),
	.rfifrdat1_9(\RF|rfif.rdat1[9]~449_combout ),
	.rfifrdat1_91(\RF|rfif.rdat1[9]~459_combout ),
	.rfifrdat2_8(\RF|rfif.rdat2[8]~503_combout ),
	.rfifrdat1_8(\RF|rfif.rdat1[8]~469_combout ),
	.rfifrdat1_81(\RF|rfif.rdat1[8]~479_combout ),
	.rfifrdat2_7(\RF|rfif.rdat2[7]~524_combout ),
	.rfifrdat1_7(\RF|rfif.rdat1[7]~489_combout ),
	.rfifrdat1_71(\RF|rfif.rdat1[7]~499_combout ),
	.rfifrdat2_6(\RF|rfif.rdat2[6]~545_combout ),
	.rfifrdat1_6(\RF|rfif.rdat1[6]~509_combout ),
	.rfifrdat1_61(\RF|rfif.rdat1[6]~519_combout ),
	.rfifrdat2_5(\RF|rfif.rdat2[5]~566_combout ),
	.rfifrdat1_5(\RF|rfif.rdat1[5]~529_combout ),
	.rfifrdat1_51(\RF|rfif.rdat1[5]~539_combout ),
	.rfifrdat2_4(\RF|rfif.rdat2[4]~587_combout ),
	.rfifrdat1_4(\RF|rfif.rdat1[4]~549_combout ),
	.rfifrdat1_41(\RF|rfif.rdat1[4]~559_combout ),
	.rfifrdat2_3(\RF|rfif.rdat2[3]~608_combout ),
	.rfifrdat1_3(\RF|rfif.rdat1[3]~569_combout ),
	.rfifrdat1_32(\RF|rfif.rdat1[3]~579_combout ),
	.rfifrdat2_2(\RF|rfif.rdat2[2]~629_combout ),
	.rfifrdat1_2(\RF|rfif.rdat1[2]~589_combout ),
	.rfifrdat1_210(\RF|rfif.rdat1[2]~599_combout ),
	.rfifrdat2_1(\RF|rfif.rdat2[1]~650_combout ),
	.rfifrdat1_1(\RF|rfif.rdat1[1]~609_combout ),
	.rfifrdat1_110(\RF|rfif.rdat1[1]~619_combout ),
	.rfifrdat2_0(\RF|rfif.rdat2[0]~671_combout ),
	.rfifrdat1_0(\RF|rfif.rdat1[0]~629_combout ),
	.rfifrdat1_01(\RF|rfif.rdat1[0]~639_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

hazard_unit HZ(
	.MemToReg_EX(MemToReg_EX),
	.RegDst_EX_0(\PR|RegDst_EX [0]),
	.RegDst_EX_1(\PR|RegDst_EX [1]),
	.RegDst_EX_2(\PR|RegDst_EX [2]),
	.RegWen_EX(\PR|RegWen_EX~q ),
	.RegDst_EX_3(\PR|RegDst_EX [3]),
	.RegDst_EX_4(\PR|RegDst_EX [4]),
	.Instr_ID_16(\PR|Instr_ID [16]),
	.hazard_Reg_ID(\PR|hazard_Reg_ID~q ),
	.Instr_ID_17(\PR|Instr_ID [17]),
	.always0(\HZ|always0~0_combout ),
	.Instr_ID_18(\PR|Instr_ID [18]),
	.Equal4(\HZ|Equal4~2_combout ),
	.Instr_ID_19(\PR|Instr_ID [19]),
	.Equal41(\HZ|Equal4~3_combout ),
	.Instr_ID_20(\PR|Instr_ID [20]),
	.Equal42(\HZ|Equal4~4_combout ),
	.MemToReg_MEM(\PR|MemToReg_MEM~q ),
	.always01(\HZ|always0~1_combout ),
	.RegWen_MEM(\PR|RegWen_MEM~q ),
	.RegDst_MEM_0(\PR|RegDst_MEM [0]),
	.output_RegWen_MEM(\output_RegWen_MEM~0_combout ),
	.RegDst_MEM_1(\PR|RegDst_MEM [1]),
	.RegDst_MEM_4(\PR|RegDst_MEM [4]),
	.output_RegWen_MEM1(\output_RegWen_MEM~1_combout ),
	.RegDst_MEM_3(\PR|RegDst_MEM [3]),
	.RegDst_MEM_2(\PR|RegDst_MEM [2]),
	.src2_hazard_t(\HZ|src2_hazard_t~2_combout ),
	.Instr_ID_21(\PR|Instr_ID [21]),
	.Instr_ID_22(\PR|Instr_ID [22]),
	.always02(\HZ|always0~2_combout ),
	.Instr_ID_24(\PR|Instr_ID [24]),
	.Equal0(\HZ|Equal0~2_combout ),
	.Instr_ID_25(\PR|Instr_ID [25]),
	.Equal01(\HZ|Equal0~3_combout ),
	.Instr_ID_23(\PR|Instr_ID [23]),
	.always03(\HZ|always0~8_combout ),
	.src1_hazard_t(\HZ|src1_hazard_t~1_combout ),
	.src2_hazard_t1(\HZ|src2_hazard_t~3_combout ),
	.src2_hazard_t2(\HZ|src2_hazard_t~4_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CU(
	.Instr_IF_30(\PR|Instr_IF [30]),
	.Instr_IF_28(\PR|Instr_IF [28]),
	.Instr_IF_26(\PR|Instr_IF [26]),
	.Instr_IF_27(\PR|Instr_IF [27]),
	.Selector14(\CU|Selector14~0_combout ),
	.Instr_IF_29(\PR|Instr_IF [29]),
	.Instr_IF_5(\PR|Instr_IF [5]),
	.Instr_IF_4(\PR|Instr_IF [4]),
	.Instr_IF_2(\PR|Instr_IF [2]),
	.Instr_IF_3(\PR|Instr_IF [3]),
	.Instr_IF_0(\PR|Instr_IF [0]),
	.Selector11(\CU|Selector11~0_combout ),
	.Instr_IF_1(\PR|Instr_IF [1]),
	.WideOr4(\CU|WideOr4~0_combout ),
	.WideOr41(\CU|WideOr4~1_combout ),
	.Instr_IF_31(\PR|Instr_IF [31]),
	.input_hazard_Reg_ID(\CU|input_hazard_Reg_ID~0_combout ),
	.WideOr21(\CU|WideOr21~0_combout ),
	.Selector141(\CU|Selector14~2_combout ),
	.WideOr211(\CU|WideOr21~2_combout ),
	.WideOr212(\CU|WideOr21~3_combout ),
	.WideOr14(\CU|WideOr14~0_combout ),
	.WideOr6(\CU|WideOr6~0_combout ),
	.WideOr61(\CU|WideOr6~1_combout ),
	.WideOr33(\CU|WideOr33~0_combout ),
	.Decoder0(\CU|Decoder0~1_combout ),
	.WideOr11(\CU|WideOr11~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline_registers PR(
	.pc_next_plus4_2(\pc_next_plus4[2]~0_combout ),
	.pc_next_plus4_3(\pc_next_plus4[3]~2_combout ),
	.pc_next_plus4_4(\pc_next_plus4[4]~4_combout ),
	.pc_next_plus4_5(\pc_next_plus4[5]~6_combout ),
	.pc_next_plus4_6(\pc_next_plus4[6]~8_combout ),
	.pc_next_plus4_7(\pc_next_plus4[7]~10_combout ),
	.pc_next_plus4_8(\pc_next_plus4[8]~12_combout ),
	.pc_next_plus4_9(\pc_next_plus4[9]~14_combout ),
	.pc_next_plus4_10(\pc_next_plus4[10]~16_combout ),
	.pc_next_plus4_11(\pc_next_plus4[11]~18_combout ),
	.pc_next_plus4_12(\pc_next_plus4[12]~20_combout ),
	.pc_next_plus4_13(\pc_next_plus4[13]~22_combout ),
	.pc_next_plus4_14(\pc_next_plus4[14]~24_combout ),
	.pc_next_plus4_15(\pc_next_plus4[15]~26_combout ),
	.pc_next_plus4_16(\pc_next_plus4[16]~28_combout ),
	.pc_next_plus4_17(\pc_next_plus4[17]~30_combout ),
	.pc_next_plus4_18(\pc_next_plus4[18]~32_combout ),
	.pc_next_plus4_19(\pc_next_plus4[19]~34_combout ),
	.pc_next_plus4_20(\pc_next_plus4[20]~36_combout ),
	.pc_next_plus4_21(\pc_next_plus4[21]~38_combout ),
	.pc_next_plus4_22(\pc_next_plus4[22]~40_combout ),
	.pc_next_plus4_23(\pc_next_plus4[23]~42_combout ),
	.pc_next_plus4_24(\pc_next_plus4[24]~44_combout ),
	.pc_next_plus4_25(\pc_next_plus4[25]~46_combout ),
	.pc_next_plus4_26(\pc_next_plus4[26]~48_combout ),
	.pc_next_plus4_27(\pc_next_plus4[27]~50_combout ),
	.pc_next_plus4_28(\pc_next_plus4[28]~52_combout ),
	.pc_next_plus4_29(\pc_next_plus4[29]~54_combout ),
	.pc_next_plus4_30(\pc_next_plus4[30]~56_combout ),
	.pc_next_plus4_31(\pc_next_plus4[31]~58_combout ),
	.Result_EX_1(Result_EX_1),
	.pc_1(pc_1),
	.Memwrite_EX1(Memwrite_EX),
	.MemToReg_EX1(MemToReg_EX),
	.Result_EX_0(Result_EX_0),
	.pc_0(pc_0),
	.Result_EX_3(Result_EX_3),
	.Result_EX_2(Result_EX_2),
	.Result_EX_5(Result_EX_5),
	.Result_EX_4(Result_EX_4),
	.Result_EX_7(Result_EX_7),
	.Result_EX_6(Result_EX_6),
	.Result_EX_9(Result_EX_9),
	.Result_EX_8(Result_EX_8),
	.Result_EX_11(Result_EX_11),
	.Result_EX_10(Result_EX_10),
	.Result_EX_13(Result_EX_13),
	.Result_EX_12(Result_EX_12),
	.Result_EX_15(Result_EX_15),
	.Result_EX_14(Result_EX_14),
	.Result_EX_17(Result_EX_17),
	.Result_EX_16(Result_EX_16),
	.Result_EX_19(Result_EX_19),
	.Result_EX_18(Result_EX_18),
	.Result_EX_21(Result_EX_21),
	.Result_EX_20(Result_EX_20),
	.Result_EX_23(Result_EX_23),
	.Result_EX_22(Result_EX_22),
	.Result_EX_25(Result_EX_25),
	.Result_EX_24(Result_EX_24),
	.Result_EX_27(Result_EX_27),
	.Result_EX_26(Result_EX_26),
	.Result_EX_29(Result_EX_29),
	.Result_EX_28(Result_EX_28),
	.Result_EX_31(Result_EX_31),
	.Result_EX_30(Result_EX_30),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.halt_MEM1(\PR|halt_MEM~q ),
	.care_ID1(\PR|care_ID~q ),
	.ALUOP_ID_1(\PR|ALUOP_ID [1]),
	.ALUOP_ID_3(\PR|ALUOP_ID [3]),
	.ALUOP_ID_2(\PR|ALUOP_ID [2]),
	.RegDst_EX_0(\PR|RegDst_EX [0]),
	.RegDst_EX_1(\PR|RegDst_EX [1]),
	.RegDst_EX_2(\PR|RegDst_EX [2]),
	.RegWen_EX1(\PR|RegWen_EX~q ),
	.RegDst_EX_3(\PR|RegDst_EX [3]),
	.RegDst_EX_4(\PR|RegDst_EX [4]),
	.Instr_ID_16(\PR|Instr_ID [16]),
	.hazard_Reg_ID1(\PR|hazard_Reg_ID~q ),
	.Instr_ID_17(\PR|Instr_ID [17]),
	.Instr_ID_18(\PR|Instr_ID [18]),
	.Instr_ID_19(\PR|Instr_ID [19]),
	.Memwrite_ID1(\PR|Memwrite_ID~q ),
	.Instr_ID_20(\PR|Instr_ID [20]),
	.ReadData_MEM_31(\PR|ReadData_MEM [31]),
	.CalcData_MEM_31(\PR|CalcData_MEM [31]),
	.MemToReg_MEM1(\PR|MemToReg_MEM~q ),
	.input_a(\input_a~56_combout ),
	.always0(\HZ|always0~1_combout ),
	.RegWen_MEM1(\PR|RegWen_MEM~q ),
	.RegDst_MEM_0(\PR|RegDst_MEM [0]),
	.RegDst_MEM_1(\PR|RegDst_MEM [1]),
	.RegDst_MEM_4(\PR|RegDst_MEM [4]),
	.RegDst_MEM_3(\PR|RegDst_MEM [3]),
	.RegDst_MEM_2(\PR|RegDst_MEM [2]),
	.ALUSrc2_ID_31(\PR|ALUSrc2_ID [31]),
	.Instr_ID_21(\PR|Instr_ID [21]),
	.Instr_ID_22(\PR|Instr_ID [22]),
	.Instr_ID_24(\PR|Instr_ID [24]),
	.Instr_ID_25(\PR|Instr_ID [25]),
	.Instr_ID_23(\PR|Instr_ID [23]),
	.ALUSrc1_ID_31(\PR|ALUSrc1_ID [31]),
	.always01(\HZ|always0~8_combout ),
	.src1_hazard_t(\HZ|src1_hazard_t~1_combout ),
	.ALUOP_ID_0(\PR|ALUOP_ID [0]),
	.ALUSrc1_ID_30(\PR|ALUSrc1_ID [30]),
	.ReadData_MEM_30(\PR|ReadData_MEM [30]),
	.CalcData_MEM_30(\PR|CalcData_MEM [30]),
	.input_b(\input_b~7_combout ),
	.ALUSrc2_ID_30(\PR|ALUSrc2_ID [30]),
	.ALUSrc1_ID_29(\PR|ALUSrc1_ID [29]),
	.ReadData_MEM_29(\PR|ReadData_MEM [29]),
	.CalcData_MEM_29(\PR|CalcData_MEM [29]),
	.input_b1(\input_b~10_combout ),
	.ALUSrc2_ID_29(\PR|ALUSrc2_ID [29]),
	.ALUSrc1_ID_28(\PR|ALUSrc1_ID [28]),
	.ReadData_MEM_28(\PR|ReadData_MEM [28]),
	.CalcData_MEM_28(\PR|CalcData_MEM [28]),
	.input_b2(\input_b~13_combout ),
	.ALUSrc2_ID_28(\PR|ALUSrc2_ID [28]),
	.ALUSrc1_ID_27(\PR|ALUSrc1_ID [27]),
	.ReadData_MEM_27(\PR|ReadData_MEM [27]),
	.CalcData_MEM_27(\PR|CalcData_MEM [27]),
	.input_b3(\input_b~16_combout ),
	.ALUSrc2_ID_27(\PR|ALUSrc2_ID [27]),
	.ALUSrc1_ID_26(\PR|ALUSrc1_ID [26]),
	.ReadData_MEM_26(\PR|ReadData_MEM [26]),
	.CalcData_MEM_26(\PR|CalcData_MEM [26]),
	.input_b4(\input_b~19_combout ),
	.ALUSrc2_ID_26(\PR|ALUSrc2_ID [26]),
	.ALUSrc1_ID_25(\PR|ALUSrc1_ID [25]),
	.ReadData_MEM_25(\PR|ReadData_MEM [25]),
	.CalcData_MEM_25(\PR|CalcData_MEM [25]),
	.input_b5(\input_b~22_combout ),
	.ALUSrc2_ID_25(\PR|ALUSrc2_ID [25]),
	.ALUSrc1_ID_24(\PR|ALUSrc1_ID [24]),
	.ReadData_MEM_24(\PR|ReadData_MEM [24]),
	.CalcData_MEM_24(\PR|CalcData_MEM [24]),
	.input_b6(\input_b~25_combout ),
	.ALUSrc2_ID_24(\PR|ALUSrc2_ID [24]),
	.ALUSrc1_ID_23(\PR|ALUSrc1_ID [23]),
	.ReadData_MEM_23(\PR|ReadData_MEM [23]),
	.CalcData_MEM_23(\PR|CalcData_MEM [23]),
	.input_b7(\input_b~28_combout ),
	.ALUSrc2_ID_23(\PR|ALUSrc2_ID [23]),
	.ALUSrc1_ID_22(\PR|ALUSrc1_ID [22]),
	.ReadData_MEM_22(\PR|ReadData_MEM [22]),
	.CalcData_MEM_22(\PR|CalcData_MEM [22]),
	.input_b8(\input_b~31_combout ),
	.ALUSrc2_ID_22(\PR|ALUSrc2_ID [22]),
	.ALUSrc1_ID_21(\PR|ALUSrc1_ID [21]),
	.ReadData_MEM_21(\PR|ReadData_MEM [21]),
	.CalcData_MEM_21(\PR|CalcData_MEM [21]),
	.input_b9(\input_b~34_combout ),
	.ALUSrc2_ID_21(\PR|ALUSrc2_ID [21]),
	.ALUSrc1_ID_20(\PR|ALUSrc1_ID [20]),
	.ReadData_MEM_20(\PR|ReadData_MEM [20]),
	.CalcData_MEM_20(\PR|CalcData_MEM [20]),
	.input_b10(\input_b~37_combout ),
	.ALUSrc2_ID_20(\PR|ALUSrc2_ID [20]),
	.ALUSrc1_ID_19(\PR|ALUSrc1_ID [19]),
	.ReadData_MEM_19(\PR|ReadData_MEM [19]),
	.CalcData_MEM_19(\PR|CalcData_MEM [19]),
	.input_b11(\input_b~40_combout ),
	.ALUSrc2_ID_19(\PR|ALUSrc2_ID [19]),
	.ALUSrc1_ID_18(\PR|ALUSrc1_ID [18]),
	.ReadData_MEM_18(\PR|ReadData_MEM [18]),
	.CalcData_MEM_18(\PR|CalcData_MEM [18]),
	.input_b12(\input_b~43_combout ),
	.ALUSrc2_ID_18(\PR|ALUSrc2_ID [18]),
	.ALUSrc1_ID_17(\PR|ALUSrc1_ID [17]),
	.ReadData_MEM_17(\PR|ReadData_MEM [17]),
	.CalcData_MEM_17(\PR|CalcData_MEM [17]),
	.input_b13(\input_b~46_combout ),
	.ALUSrc2_ID_17(\PR|ALUSrc2_ID [17]),
	.ALUSrc1_ID_16(\PR|ALUSrc1_ID [16]),
	.ReadData_MEM_16(\PR|ReadData_MEM [16]),
	.CalcData_MEM_16(\PR|CalcData_MEM [16]),
	.input_b14(\input_b~49_combout ),
	.ALUSrc2_ID_16(\PR|ALUSrc2_ID [16]),
	.ALUSrc1_ID_15(\PR|ALUSrc1_ID [15]),
	.ReadData_MEM_15(\PR|ReadData_MEM [15]),
	.CalcData_MEM_15(\PR|CalcData_MEM [15]),
	.input_b15(\input_b~52_combout ),
	.ALUSrc2_ID_15(\PR|ALUSrc2_ID [15]),
	.ALUSrc1_ID_14(\PR|ALUSrc1_ID [14]),
	.ReadData_MEM_14(\PR|ReadData_MEM [14]),
	.CalcData_MEM_14(\PR|CalcData_MEM [14]),
	.input_b16(\input_b~55_combout ),
	.ALUSrc2_ID_14(\PR|ALUSrc2_ID [14]),
	.ReadData_MEM_13(\PR|ReadData_MEM [13]),
	.CalcData_MEM_13(\PR|CalcData_MEM [13]),
	.input_a1(\input_a~96_combout ),
	.ALUSrc2_ID_13(\PR|ALUSrc2_ID [13]),
	.ALUSrc1_ID_13(\PR|ALUSrc1_ID [13]),
	.ReadData_MEM_12(\PR|ReadData_MEM [12]),
	.CalcData_MEM_12(\PR|CalcData_MEM [12]),
	.input_a2(\input_a~99_combout ),
	.ALUSrc2_ID_12(\PR|ALUSrc2_ID [12]),
	.ALUSrc1_ID_12(\PR|ALUSrc1_ID [12]),
	.ReadData_MEM_11(\PR|ReadData_MEM [11]),
	.CalcData_MEM_11(\PR|CalcData_MEM [11]),
	.input_a3(\input_a~102_combout ),
	.ALUSrc2_ID_11(\PR|ALUSrc2_ID [11]),
	.ALUSrc1_ID_11(\PR|ALUSrc1_ID [11]),
	.ReadData_MEM_10(\PR|ReadData_MEM [10]),
	.CalcData_MEM_10(\PR|CalcData_MEM [10]),
	.input_a4(\input_a~105_combout ),
	.ALUSrc2_ID_10(\PR|ALUSrc2_ID [10]),
	.ALUSrc1_ID_10(\PR|ALUSrc1_ID [10]),
	.ReadData_MEM_9(\PR|ReadData_MEM [9]),
	.CalcData_MEM_9(\PR|CalcData_MEM [9]),
	.input_a5(\input_a~108_combout ),
	.ALUSrc2_ID_9(\PR|ALUSrc2_ID [9]),
	.ALUSrc1_ID_9(\PR|ALUSrc1_ID [9]),
	.ReadData_MEM_8(\PR|ReadData_MEM [8]),
	.CalcData_MEM_8(\PR|CalcData_MEM [8]),
	.input_a6(\input_a~111_combout ),
	.ALUSrc2_ID_8(\PR|ALUSrc2_ID [8]),
	.ALUSrc1_ID_8(\PR|ALUSrc1_ID [8]),
	.ReadData_MEM_7(\PR|ReadData_MEM [7]),
	.CalcData_MEM_7(\PR|CalcData_MEM [7]),
	.input_a7(\input_a~114_combout ),
	.ALUSrc2_ID_7(\PR|ALUSrc2_ID [7]),
	.ALUSrc1_ID_7(\PR|ALUSrc1_ID [7]),
	.ReadData_MEM_6(\PR|ReadData_MEM [6]),
	.CalcData_MEM_6(\PR|CalcData_MEM [6]),
	.input_a8(\input_a~117_combout ),
	.ALUSrc2_ID_6(\PR|ALUSrc2_ID [6]),
	.ALUSrc1_ID_6(\PR|ALUSrc1_ID [6]),
	.ReadData_MEM_5(\PR|ReadData_MEM [5]),
	.CalcData_MEM_5(\PR|CalcData_MEM [5]),
	.input_a9(\input_a~120_combout ),
	.ALUSrc2_ID_5(\PR|ALUSrc2_ID [5]),
	.ALUSrc1_ID_5(\PR|ALUSrc1_ID [5]),
	.ReadData_MEM_4(\PR|ReadData_MEM [4]),
	.CalcData_MEM_4(\PR|CalcData_MEM [4]),
	.input_a10(\input_a~123_combout ),
	.ALUSrc2_ID_4(\PR|ALUSrc2_ID [4]),
	.ALUSrc1_ID_4(\PR|ALUSrc1_ID [4]),
	.ReadData_MEM_3(\PR|ReadData_MEM [3]),
	.CalcData_MEM_3(\PR|CalcData_MEM [3]),
	.input_a11(\input_a~126_combout ),
	.ALUSrc2_ID_3(\PR|ALUSrc2_ID [3]),
	.ALUSrc1_ID_3(\PR|ALUSrc1_ID [3]),
	.ReadData_MEM_2(\PR|ReadData_MEM [2]),
	.CalcData_MEM_2(\PR|CalcData_MEM [2]),
	.input_a12(\input_a~129_combout ),
	.ALUSrc2_ID_2(\PR|ALUSrc2_ID [2]),
	.ALUSrc1_ID_2(\PR|ALUSrc1_ID [2]),
	.ReadData_MEM_1(\PR|ReadData_MEM [1]),
	.CalcData_MEM_1(\PR|CalcData_MEM [1]),
	.input_a13(\input_a~132_combout ),
	.ALUSrc2_ID_1(\PR|ALUSrc2_ID [1]),
	.ALUSrc1_ID_1(\PR|ALUSrc1_ID [1]),
	.ReadData_MEM_0(\PR|ReadData_MEM [0]),
	.CalcData_MEM_0(\PR|CalcData_MEM [0]),
	.input_a14(\input_a~135_combout ),
	.ALUSrc2_ID_0(\PR|ALUSrc2_ID [0]),
	.ALUSrc1_ID_0(\PR|ALUSrc1_ID [0]),
	.Wdata_EX_0(Wdata_EX_0),
	.src2_hazard_t(\HZ|src2_hazard_t~3_combout ),
	.nextPC_ID_1(\PR|nextPC_ID [1]),
	.Selector30(\ALU|Selector30~7_combout ),
	.jump_ID_0(\PR|jump_ID [0]),
	.jump_ID_1(\PR|jump_ID [1]),
	.jump_ID_2(\PR|jump_ID [2]),
	.Equal8(\Equal8~0_combout ),
	.Selector28(\ALU|Selector28~10_combout ),
	.Selector3(\ALU|Selector3~11_combout ),
	.Selector22(\ALU|Selector22~9_combout ),
	.Selector2(\ALU|Selector2~8_combout ),
	.Selector27(\ALU|Selector27~8_combout ),
	.Selector25(\ALU|Selector25~7_combout ),
	.Selector24(\ALU|Selector24~8_combout ),
	.Selector26(\ALU|Selector26~7_combout ),
	.Selector4(\ALU|Selector4~7_combout ),
	.Selector16(\ALU|Selector16~10_combout ),
	.Selector7(\ALU|Selector7~12_combout ),
	.Selector6(\ALU|Selector6~6_combout ),
	.Selector29(\ALU|Selector29~10_combout ),
	.Selector15(\ALU|Selector15~14_combout ),
	.Selector5(\ALU|Selector5~6_combout ),
	.Selector31(\ALU|Selector31~11_combout ),
	.Selector11(\ALU|Selector11~9_combout ),
	.Selector10(\ALU|Selector10~8_combout ),
	.Selector21(\ALU|Selector21~9_combout ),
	.Selector20(\ALU|Selector20~8_combout ),
	.Selector9(\ALU|Selector9~8_combout ),
	.Selector8(\ALU|Selector8~8_combout ),
	.Selector14(\ALU|Selector14~7_combout ),
	.Selector13(\ALU|Selector13~7_combout ),
	.Selector12(\ALU|Selector12~7_combout ),
	.Selector23(\ALU|Selector23~10_combout ),
	.Selector19(\ALU|Selector19~9_combout ),
	.Selector18(\ALU|Selector18~8_combout ),
	.Selector17(\ALU|Selector17~7_combout ),
	.Selector0(\ALU|Selector0~28_combout ),
	.Selector1(\ALU|Selector1~11_combout ),
	.branch(\branch~0_combout ),
	.always02(always0),
	.nextPC_ID_0(\PR|nextPC_ID [0]),
	.nextPC_ID_3(\PR|nextPC_ID [3]),
	.Instr_ID_1(\PR|Instr_ID [1]),
	.nextPC_ID_2(\PR|nextPC_ID [2]),
	.Instr_ID_0(\PR|Instr_ID [0]),
	.nextPC_ID_5(\PR|nextPC_ID [5]),
	.Instr_ID_3(\PR|Instr_ID [3]),
	.nextPC_ID_4(\PR|nextPC_ID [4]),
	.Instr_ID_2(\PR|Instr_ID [2]),
	.nextPC_ID_7(\PR|nextPC_ID [7]),
	.Instr_ID_5(\PR|Instr_ID [5]),
	.nextPC_ID_6(\PR|nextPC_ID [6]),
	.Instr_ID_4(\PR|Instr_ID [4]),
	.nextPC_ID_9(\PR|nextPC_ID [9]),
	.Instr_ID_7(\PR|Instr_ID [7]),
	.nextPC_ID_8(\PR|nextPC_ID [8]),
	.Instr_ID_6(\PR|Instr_ID [6]),
	.nextPC_ID_11(\PR|nextPC_ID [11]),
	.Instr_ID_9(\PR|Instr_ID [9]),
	.nextPC_ID_10(\PR|nextPC_ID [10]),
	.Instr_ID_8(\PR|Instr_ID [8]),
	.nextPC_ID_13(\PR|nextPC_ID [13]),
	.Instr_ID_11(\PR|Instr_ID [11]),
	.nextPC_ID_12(\PR|nextPC_ID [12]),
	.Instr_ID_10(\PR|Instr_ID [10]),
	.nextPC_ID_15(\PR|nextPC_ID [15]),
	.Instr_ID_13(\PR|Instr_ID [13]),
	.nextPC_ID_14(\PR|nextPC_ID [14]),
	.Instr_ID_12(\PR|Instr_ID [12]),
	.nextPC_ID_17(\PR|nextPC_ID [17]),
	.Instr_ID_15(\PR|Instr_ID [15]),
	.nextPC_ID_16(\PR|nextPC_ID [16]),
	.Instr_ID_14(\PR|Instr_ID [14]),
	.nextPC_ID_19(\PR|nextPC_ID [19]),
	.nextPC_ID_18(\PR|nextPC_ID [18]),
	.nextPC_ID_21(\PR|nextPC_ID [21]),
	.nextPC_ID_20(\PR|nextPC_ID [20]),
	.nextPC_ID_23(\PR|nextPC_ID [23]),
	.nextPC_ID_22(\PR|nextPC_ID [22]),
	.nextPC_ID_25(\PR|nextPC_ID [25]),
	.nextPC_ID_24(\PR|nextPC_ID [24]),
	.nextPC_ID_27(\PR|nextPC_ID [27]),
	.nextPC_ID_26(\PR|nextPC_ID [26]),
	.nextPC_ID_29(\PR|nextPC_ID [29]),
	.nextPC_ID_28(\PR|nextPC_ID [28]),
	.nextPC_ID_31(\PR|nextPC_ID [31]),
	.nextPC_ID_30(\PR|nextPC_ID [30]),
	.Wdata_EX_1(Wdata_EX_1),
	.Wdata_EX_2(Wdata_EX_2),
	.Wdata_EX_3(Wdata_EX_3),
	.Wdata_EX_4(Wdata_EX_4),
	.Wdata_EX_5(Wdata_EX_5),
	.Wdata_EX_6(Wdata_EX_6),
	.Wdata_EX_7(Wdata_EX_7),
	.Wdata_EX_8(Wdata_EX_8),
	.Wdata_EX_9(Wdata_EX_9),
	.Wdata_EX_10(Wdata_EX_10),
	.Wdata_EX_11(Wdata_EX_11),
	.Wdata_EX_12(Wdata_EX_12),
	.Wdata_EX_13(Wdata_EX_13),
	.Wdata_EX_14(Wdata_EX_14),
	.Wdata_EX_15(Wdata_EX_15),
	.Wdata_EX_16(Wdata_EX_16),
	.Wdata_EX_17(Wdata_EX_17),
	.Wdata_EX_18(Wdata_EX_18),
	.Wdata_EX_19(Wdata_EX_19),
	.Wdata_EX_20(Wdata_EX_20),
	.Wdata_EX_21(Wdata_EX_21),
	.Wdata_EX_22(Wdata_EX_22),
	.Wdata_EX_23(Wdata_EX_23),
	.Wdata_EX_24(Wdata_EX_24),
	.Wdata_EX_25(Wdata_EX_25),
	.Wdata_EX_26(Wdata_EX_26),
	.Wdata_EX_27(Wdata_EX_27),
	.Wdata_EX_28(Wdata_EX_28),
	.Wdata_EX_29(Wdata_EX_29),
	.Wdata_EX_30(Wdata_EX_30),
	.Wdata_EX_31(Wdata_EX_31),
	.Instr_IF_30(\PR|Instr_IF [30]),
	.Instr_IF_28(\PR|Instr_IF [28]),
	.Instr_IF_26(\PR|Instr_IF [26]),
	.Instr_IF_27(\PR|Instr_IF [27]),
	.Selector141(\CU|Selector14~0_combout ),
	.Instr_IF_29(\PR|Instr_IF [29]),
	.Instr_IF_5(\PR|Instr_IF [5]),
	.Instr_IF_4(\PR|Instr_IF [4]),
	.Instr_IF_2(\PR|Instr_IF [2]),
	.Instr_IF_3(\PR|Instr_IF [3]),
	.Instr_IF_0(\PR|Instr_IF [0]),
	.src2_hazard_t1(\HZ|src2_hazard_t~4_combout ),
	.Selector111(\CU|Selector11~0_combout ),
	.Instr_IF_1(\PR|Instr_IF [1]),
	.WideOr4(\CU|WideOr4~0_combout ),
	.WideOr41(\CU|WideOr4~1_combout ),
	.Instr_IF_31(\PR|Instr_IF [31]),
	.Instr_IF_16(\PR|Instr_IF [16]),
	.input_hazard_Reg_ID(\CU|input_hazard_Reg_ID~0_combout ),
	.Instr_IF_17(\PR|Instr_IF [17]),
	.Instr_IF_18(\PR|Instr_IF [18]),
	.Instr_IF_19(\PR|Instr_IF [19]),
	.WideOr21(\CU|WideOr21~0_combout ),
	.Instr_IF_20(\PR|Instr_IF [20]),
	.Equal20(\Equal20~0_combout ),
	.Selector142(\CU|Selector14~2_combout ),
	.WideOr211(\CU|WideOr21~2_combout ),
	.WideOr212(\CU|WideOr21~3_combout ),
	.rfifrdat2_31(\RF|rfif.rdat2[31]~20_combout ),
	.WideOr14(\CU|WideOr14~0_combout ),
	.Instr_IF_21(\PR|Instr_IF [21]),
	.Instr_IF_22(\PR|Instr_IF [22]),
	.Instr_IF_24(\PR|Instr_IF [24]),
	.Instr_IF_25(\PR|Instr_IF [25]),
	.Instr_IF_23(\PR|Instr_IF [23]),
	.rfifrdat1_31(\RF|rfif.rdat1[31]~9_combout ),
	.rfifrdat1_311(\RF|rfif.rdat1[31]~19_combout ),
	.WideOr0(\RF|WideOr0~0_combout ),
	.WideOr6(\CU|WideOr6~0_combout ),
	.WideOr61(\CU|WideOr6~1_combout ),
	.rfifrdat1_30(\RF|rfif.rdat1[30]~29_combout ),
	.rfifrdat1_301(\RF|rfif.rdat1[30]~39_combout ),
	.rfifrdat2_30(\RF|rfif.rdat2[30]~41_combout ),
	.rfifrdat1_29(\RF|rfif.rdat1[29]~49_combout ),
	.rfifrdat1_291(\RF|rfif.rdat1[29]~59_combout ),
	.rfifrdat2_29(\RF|rfif.rdat2[29]~62_combout ),
	.rfifrdat1_28(\RF|rfif.rdat1[28]~69_combout ),
	.rfifrdat1_281(\RF|rfif.rdat1[28]~79_combout ),
	.rfifrdat2_28(\RF|rfif.rdat2[28]~83_combout ),
	.rfifrdat1_27(\RF|rfif.rdat1[27]~89_combout ),
	.rfifrdat1_271(\RF|rfif.rdat1[27]~99_combout ),
	.rfifrdat2_27(\RF|rfif.rdat2[27]~104_combout ),
	.rfifrdat1_26(\RF|rfif.rdat1[26]~109_combout ),
	.rfifrdat1_261(\RF|rfif.rdat1[26]~119_combout ),
	.rfifrdat2_26(\RF|rfif.rdat2[26]~125_combout ),
	.Instr_IF_10(\PR|Instr_IF [10]),
	.rfifrdat1_25(\RF|rfif.rdat1[25]~129_combout ),
	.rfifrdat1_251(\RF|rfif.rdat1[25]~139_combout ),
	.rfifrdat2_25(\RF|rfif.rdat2[25]~146_combout ),
	.Instr_IF_9(\PR|Instr_IF [9]),
	.rfifrdat1_24(\RF|rfif.rdat1[24]~149_combout ),
	.rfifrdat1_241(\RF|rfif.rdat1[24]~159_combout ),
	.rfifrdat2_24(\RF|rfif.rdat2[24]~167_combout ),
	.Instr_IF_8(\PR|Instr_IF [8]),
	.rfifrdat1_23(\RF|rfif.rdat1[23]~169_combout ),
	.rfifrdat1_231(\RF|rfif.rdat1[23]~179_combout ),
	.rfifrdat2_23(\RF|rfif.rdat2[23]~188_combout ),
	.Instr_IF_7(\PR|Instr_IF [7]),
	.rfifrdat1_22(\RF|rfif.rdat1[22]~189_combout ),
	.rfifrdat1_221(\RF|rfif.rdat1[22]~199_combout ),
	.rfifrdat2_22(\RF|rfif.rdat2[22]~209_combout ),
	.Instr_IF_6(\PR|Instr_IF [6]),
	.rfifrdat1_21(\RF|rfif.rdat1[21]~209_combout ),
	.rfifrdat1_211(\RF|rfif.rdat1[21]~219_combout ),
	.rfifrdat2_21(\RF|rfif.rdat2[21]~230_combout ),
	.rfifrdat1_20(\RF|rfif.rdat1[20]~229_combout ),
	.rfifrdat1_201(\RF|rfif.rdat1[20]~239_combout ),
	.rfifrdat2_20(\RF|rfif.rdat2[20]~251_combout ),
	.rfifrdat1_19(\RF|rfif.rdat1[19]~249_combout ),
	.rfifrdat1_191(\RF|rfif.rdat1[19]~259_combout ),
	.rfifrdat2_19(\RF|rfif.rdat2[19]~272_combout ),
	.rfifrdat1_18(\RF|rfif.rdat1[18]~269_combout ),
	.rfifrdat1_181(\RF|rfif.rdat1[18]~279_combout ),
	.rfifrdat2_18(\RF|rfif.rdat2[18]~293_combout ),
	.rfifrdat1_17(\RF|rfif.rdat1[17]~289_combout ),
	.rfifrdat1_171(\RF|rfif.rdat1[17]~299_combout ),
	.rfifrdat2_17(\RF|rfif.rdat2[17]~314_combout ),
	.rfifrdat1_16(\RF|rfif.rdat1[16]~309_combout ),
	.rfifrdat1_161(\RF|rfif.rdat1[16]~319_combout ),
	.rfifrdat2_16(\RF|rfif.rdat2[16]~335_combout ),
	.rfifrdat1_15(\RF|rfif.rdat1[15]~329_combout ),
	.rfifrdat1_151(\RF|rfif.rdat1[15]~339_combout ),
	.Equal0(\Equal0~0_combout ),
	.rfifrdat2_15(\RF|rfif.rdat2[15]~356_combout ),
	.rfifrdat1_14(\RF|rfif.rdat1[14]~349_combout ),
	.rfifrdat1_141(\RF|rfif.rdat1[14]~359_combout ),
	.rfifrdat2_14(\RF|rfif.rdat2[14]~377_combout ),
	.rfifrdat2_13(\RF|rfif.rdat2[13]~398_combout ),
	.rfifrdat1_13(\RF|rfif.rdat1[13]~369_combout ),
	.rfifrdat1_131(\RF|rfif.rdat1[13]~379_combout ),
	.rfifrdat2_12(\RF|rfif.rdat2[12]~419_combout ),
	.rfifrdat1_12(\RF|rfif.rdat1[12]~389_combout ),
	.rfifrdat1_121(\RF|rfif.rdat1[12]~399_combout ),
	.rfifrdat2_11(\RF|rfif.rdat2[11]~440_combout ),
	.rfifrdat1_11(\RF|rfif.rdat1[11]~409_combout ),
	.rfifrdat1_111(\RF|rfif.rdat1[11]~419_combout ),
	.rfifrdat2_10(\RF|rfif.rdat2[10]~461_combout ),
	.rfifrdat1_10(\RF|rfif.rdat1[10]~429_combout ),
	.rfifrdat1_101(\RF|rfif.rdat1[10]~439_combout ),
	.rfifrdat2_9(\RF|rfif.rdat2[9]~482_combout ),
	.rfifrdat1_9(\RF|rfif.rdat1[9]~449_combout ),
	.rfifrdat1_91(\RF|rfif.rdat1[9]~459_combout ),
	.rfifrdat2_8(\RF|rfif.rdat2[8]~503_combout ),
	.rfifrdat1_8(\RF|rfif.rdat1[8]~469_combout ),
	.rfifrdat1_81(\RF|rfif.rdat1[8]~479_combout ),
	.rfifrdat2_7(\RF|rfif.rdat2[7]~524_combout ),
	.rfifrdat1_7(\RF|rfif.rdat1[7]~489_combout ),
	.rfifrdat1_71(\RF|rfif.rdat1[7]~499_combout ),
	.rfifrdat2_6(\RF|rfif.rdat2[6]~545_combout ),
	.rfifrdat1_6(\RF|rfif.rdat1[6]~509_combout ),
	.rfifrdat1_61(\RF|rfif.rdat1[6]~519_combout ),
	.rfifrdat2_5(\RF|rfif.rdat2[5]~566_combout ),
	.rfifrdat1_5(\RF|rfif.rdat1[5]~529_combout ),
	.rfifrdat1_51(\RF|rfif.rdat1[5]~539_combout ),
	.rfifrdat2_4(\RF|rfif.rdat2[4]~587_combout ),
	.input_ALUSrc2_ID(\input_ALUSrc2_ID~3_combout ),
	.rfifrdat1_4(\RF|rfif.rdat1[4]~549_combout ),
	.rfifrdat1_41(\RF|rfif.rdat1[4]~559_combout ),
	.rfifrdat2_3(\RF|rfif.rdat2[3]~608_combout ),
	.input_ALUSrc2_ID1(\input_ALUSrc2_ID~5_combout ),
	.rfifrdat1_3(\RF|rfif.rdat1[3]~569_combout ),
	.rfifrdat1_32(\RF|rfif.rdat1[3]~579_combout ),
	.rfifrdat2_2(\RF|rfif.rdat2[2]~629_combout ),
	.input_ALUSrc2_ID2(\input_ALUSrc2_ID~7_combout ),
	.rfifrdat1_2(\RF|rfif.rdat1[2]~589_combout ),
	.rfifrdat1_210(\RF|rfif.rdat1[2]~599_combout ),
	.rfifrdat2_1(\RF|rfif.rdat2[1]~650_combout ),
	.input_ALUSrc2_ID3(\input_ALUSrc2_ID~9_combout ),
	.rfifrdat1_1(\RF|rfif.rdat1[1]~609_combout ),
	.rfifrdat1_110(\RF|rfif.rdat1[1]~619_combout ),
	.rfifrdat2_0(\RF|rfif.rdat2[0]~671_combout ),
	.input_ALUSrc2_ID4(\input_ALUSrc2_ID~11_combout ),
	.rfifrdat1_0(\RF|rfif.rdat1[0]~629_combout ),
	.rfifrdat1_01(\RF|rfif.rdat1[0]~639_combout ),
	.Equal27(\Equal27~0_combout ),
	.WideOr33(\CU|WideOr33~0_combout ),
	.Decoder0(\CU|Decoder0~1_combout ),
	.WideOr11(\CU|WideOr11~0_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu_file ALU(
	.Add1(\ALU|Add1~62_combout ),
	.Add0(\ALU|Add0~42_combout ),
	.Add01(\ALU|Add0~44_combout ),
	.Add02(\ALU|Add0~46_combout ),
	.Add03(\ALU|Add0~48_combout ),
	.Add04(\ALU|Add0~50_combout ),
	.Add05(\ALU|Add0~52_combout ),
	.Add06(\ALU|Add0~54_combout ),
	.Add07(\ALU|Add0~56_combout ),
	.Add08(\ALU|Add0~58_combout ),
	.Add09(\ALU|Add0~60_combout ),
	.Add010(\ALU|Add0~62_combout ),
	.Result_EX_1(Result_EX_1),
	.Result_EX_0(Result_EX_0),
	.Result_EX_3(Result_EX_3),
	.Result_EX_2(Result_EX_2),
	.Result_EX_4(Result_EX_4),
	.Result_EX_7(Result_EX_7),
	.Result_EX_31(Result_EX_31),
	.ALUOP_ID_1(\PR|ALUOP_ID [1]),
	.ALUOP_ID_3(\PR|ALUOP_ID [3]),
	.ALUOP_ID_2(\PR|ALUOP_ID [2]),
	.input_b(\input_b~1_combout ),
	.input_b1(\input_b~5_combout ),
	.input_a(\input_a~61_combout ),
	.out(\ALU|out~0_combout ),
	.ALUOP_ID_0(\PR|ALUOP_ID [0]),
	.input_b2(\input_b~6_combout ),
	.input_a1(\input_a~63_combout ),
	.input_b3(\input_b~9_combout ),
	.input_a2(\input_a~65_combout ),
	.input_b4(\input_b~12_combout ),
	.input_a3(\input_a~67_combout ),
	.input_b5(\input_b~15_combout ),
	.input_a4(\input_a~69_combout ),
	.input_b6(\input_b~18_combout ),
	.input_a5(\input_a~71_combout ),
	.input_b7(\input_b~21_combout ),
	.input_a6(\input_a~73_combout ),
	.input_b8(\input_b~24_combout ),
	.input_a7(\input_a~75_combout ),
	.input_b9(\input_b~27_combout ),
	.input_a8(\input_a~77_combout ),
	.input_b10(\input_b~30_combout ),
	.input_a9(\input_a~79_combout ),
	.input_b11(\input_b~33_combout ),
	.input_a10(\input_a~81_combout ),
	.input_b12(\input_b~36_combout ),
	.input_a11(\input_a~83_combout ),
	.input_b13(\input_b~39_combout ),
	.input_a12(\input_a~85_combout ),
	.input_b14(\input_b~42_combout ),
	.input_a13(\input_a~87_combout ),
	.input_b15(\input_b~45_combout ),
	.input_a14(\input_a~89_combout ),
	.input_b16(\input_b~48_combout ),
	.input_a15(\input_a~91_combout ),
	.input_b17(\input_b~51_combout ),
	.input_a16(\input_a~93_combout ),
	.input_b18(\input_b~54_combout ),
	.input_a17(\input_a~95_combout ),
	.input_b19(\input_b~57_combout ),
	.input_b20(\input_b~59_combout ),
	.input_a18(\input_a~98_combout ),
	.input_b21(\input_b~61_combout ),
	.input_a19(\input_a~101_combout ),
	.input_b22(\input_b~63_combout ),
	.input_a20(\input_a~104_combout ),
	.input_b23(\input_b~65_combout ),
	.input_a21(\input_a~107_combout ),
	.input_b24(\input_b~67_combout ),
	.input_a22(\input_a~110_combout ),
	.input_b25(\input_b~69_combout ),
	.input_a23(\input_a~113_combout ),
	.input_b26(\input_b~70_combout ),
	.input_b27(\input_b~71_combout ),
	.input_a24(\input_a~116_combout ),
	.input_b28(\input_b~73_combout ),
	.input_a25(\input_a~119_combout ),
	.input_b29(\input_b~75_combout ),
	.input_a26(\input_a~122_combout ),
	.input_b30(\input_b~76_combout ),
	.input_b31(\input_b~77_combout ),
	.input_a27(\input_a~125_combout ),
	.input_b32(\input_b~78_combout ),
	.input_b33(\input_b~79_combout ),
	.input_a28(\input_a~128_combout ),
	.input_b34(\input_b~80_combout ),
	.input_b35(\input_b~81_combout ),
	.input_a29(\input_a~131_combout ),
	.input_b36(\input_b~82_combout ),
	.input_b37(\input_b~83_combout ),
	.input_a30(\input_a~134_combout ),
	.input_b38(\input_b~84_combout ),
	.input_b39(\input_b~85_combout ),
	.input_a31(\input_a~137_combout ),
	.Equal0(\ALU|Equal0~0_combout ),
	.Equal01(\ALU|Equal0~5_combout ),
	.Equal02(\ALU|Equal0~6_combout ),
	.Selector30(\ALU|Selector30~7_combout ),
	.halt_reg(\halt_reg~10_combout ),
	.Selector28(\ALU|Selector28~10_combout ),
	.Selector3(\ALU|Selector3~11_combout ),
	.Selector22(\ALU|Selector22~9_combout ),
	.Selector2(\ALU|Selector2~8_combout ),
	.Selector27(\ALU|Selector27~8_combout ),
	.Selector25(\ALU|Selector25~7_combout ),
	.input_b40(\input_b~86_combout ),
	.Selector24(\ALU|Selector24~8_combout ),
	.Selector26(\ALU|Selector26~7_combout ),
	.Selector4(\ALU|Selector4~7_combout ),
	.Selector16(\ALU|Selector16~10_combout ),
	.Selector7(\ALU|Selector7~12_combout ),
	.Selector6(\ALU|Selector6~6_combout ),
	.Selector29(\ALU|Selector29~10_combout ),
	.Selector15(\ALU|Selector15~14_combout ),
	.Selector5(\ALU|Selector5~6_combout ),
	.Selector31(\ALU|Selector31~11_combout ),
	.Selector11(\ALU|Selector11~9_combout ),
	.Selector10(\ALU|Selector10~8_combout ),
	.Selector21(\ALU|Selector21~9_combout ),
	.Selector20(\ALU|Selector20~8_combout ),
	.Selector9(\ALU|Selector9~8_combout ),
	.Selector8(\ALU|Selector8~8_combout ),
	.Selector14(\ALU|Selector14~7_combout ),
	.Selector13(\ALU|Selector13~7_combout ),
	.Selector12(\ALU|Selector12~7_combout ),
	.Selector23(\ALU|Selector23~10_combout ),
	.Selector19(\ALU|Selector19~9_combout ),
	.Selector18(\ALU|Selector18~8_combout ),
	.Selector17(\ALU|Selector17~7_combout ),
	.Selector0(\ALU|Selector0~28_combout ),
	.Selector1(\ALU|Selector1~11_combout ),
	.Equal11(\ALU|Equal11~11_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \pc_next_branch[2]~0 (
// Equation(s):
// \pc_next_branch[2]~0_combout  = (nextPC_ID_2 & (Instr_ID_0 $ (VCC))) # (!nextPC_ID_2 & (Instr_ID_0 & VCC))
// \pc_next_branch[2]~1  = CARRY((nextPC_ID_2 & Instr_ID_0))

	.dataa(\PR|nextPC_ID [2]),
	.datab(\PR|Instr_ID [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pc_next_branch[2]~0_combout ),
	.cout(\pc_next_branch[2]~1 ));
// synopsys translate_off
defparam \pc_next_branch[2]~0 .lut_mask = 16'h6688;
defparam \pc_next_branch[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \pc_next_branch[8]~12 (
// Equation(s):
// \pc_next_branch[8]~12_combout  = ((nextPC_ID_8 $ (Instr_ID_6 $ (!\pc_next_branch[7]~11 )))) # (GND)
// \pc_next_branch[8]~13  = CARRY((nextPC_ID_8 & ((Instr_ID_6) # (!\pc_next_branch[7]~11 ))) # (!nextPC_ID_8 & (Instr_ID_6 & !\pc_next_branch[7]~11 )))

	.dataa(\PR|nextPC_ID [8]),
	.datab(\PR|Instr_ID [6]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[7]~11 ),
	.combout(\pc_next_branch[8]~12_combout ),
	.cout(\pc_next_branch[8]~13 ));
// synopsys translate_off
defparam \pc_next_branch[8]~12 .lut_mask = 16'h698E;
defparam \pc_next_branch[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \pc_next_branch[16]~28 (
// Equation(s):
// \pc_next_branch[16]~28_combout  = ((nextPC_ID_16 $ (Instr_ID_14 $ (!\pc_next_branch[15]~27 )))) # (GND)
// \pc_next_branch[16]~29  = CARRY((nextPC_ID_16 & ((Instr_ID_14) # (!\pc_next_branch[15]~27 ))) # (!nextPC_ID_16 & (Instr_ID_14 & !\pc_next_branch[15]~27 )))

	.dataa(\PR|nextPC_ID [16]),
	.datab(\PR|Instr_ID [14]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[15]~27 ),
	.combout(\pc_next_branch[16]~28_combout ),
	.cout(\pc_next_branch[16]~29 ));
// synopsys translate_off
defparam \pc_next_branch[16]~28 .lut_mask = 16'h698E;
defparam \pc_next_branch[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N0
cycloneive_lcell_comb \pc_next_branch[17]~30 (
// Equation(s):
// \pc_next_branch[17]~30_combout  = (nextPC_ID_17 & ((Instr_ID_15 & (\pc_next_branch[16]~29  & VCC)) # (!Instr_ID_15 & (!\pc_next_branch[16]~29 )))) # (!nextPC_ID_17 & ((Instr_ID_15 & (!\pc_next_branch[16]~29 )) # (!Instr_ID_15 & ((\pc_next_branch[16]~29 ) 
// # (GND)))))
// \pc_next_branch[17]~31  = CARRY((nextPC_ID_17 & (!Instr_ID_15 & !\pc_next_branch[16]~29 )) # (!nextPC_ID_17 & ((!\pc_next_branch[16]~29 ) # (!Instr_ID_15))))

	.dataa(\PR|nextPC_ID [17]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[16]~29 ),
	.combout(\pc_next_branch[17]~30_combout ),
	.cout(\pc_next_branch[17]~31 ));
// synopsys translate_off
defparam \pc_next_branch[17]~30 .lut_mask = 16'h9617;
defparam \pc_next_branch[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N2
cycloneive_lcell_comb \pc_next_branch[18]~32 (
// Equation(s):
// \pc_next_branch[18]~32_combout  = ((nextPC_ID_18 $ (Instr_ID_15 $ (!\pc_next_branch[17]~31 )))) # (GND)
// \pc_next_branch[18]~33  = CARRY((nextPC_ID_18 & ((Instr_ID_15) # (!\pc_next_branch[17]~31 ))) # (!nextPC_ID_18 & (Instr_ID_15 & !\pc_next_branch[17]~31 )))

	.dataa(\PR|nextPC_ID [18]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[17]~31 ),
	.combout(\pc_next_branch[18]~32_combout ),
	.cout(\pc_next_branch[18]~33 ));
// synopsys translate_off
defparam \pc_next_branch[18]~32 .lut_mask = 16'h698E;
defparam \pc_next_branch[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \pc_next_branch[20]~36 (
// Equation(s):
// \pc_next_branch[20]~36_combout  = ((nextPC_ID_20 $ (Instr_ID_15 $ (!\pc_next_branch[19]~35 )))) # (GND)
// \pc_next_branch[20]~37  = CARRY((nextPC_ID_20 & ((Instr_ID_15) # (!\pc_next_branch[19]~35 ))) # (!nextPC_ID_20 & (Instr_ID_15 & !\pc_next_branch[19]~35 )))

	.dataa(\PR|nextPC_ID [20]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[19]~35 ),
	.combout(\pc_next_branch[20]~36_combout ),
	.cout(\pc_next_branch[20]~37 ));
// synopsys translate_off
defparam \pc_next_branch[20]~36 .lut_mask = 16'h698E;
defparam \pc_next_branch[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N24
cycloneive_lcell_comb \pc_next_branch[29]~54 (
// Equation(s):
// \pc_next_branch[29]~54_combout  = (Instr_ID_15 & ((nextPC_ID_29 & (\pc_next_branch[28]~53  & VCC)) # (!nextPC_ID_29 & (!\pc_next_branch[28]~53 )))) # (!Instr_ID_15 & ((nextPC_ID_29 & (!\pc_next_branch[28]~53 )) # (!nextPC_ID_29 & ((\pc_next_branch[28]~53 
// ) # (GND)))))
// \pc_next_branch[29]~55  = CARRY((Instr_ID_15 & (!nextPC_ID_29 & !\pc_next_branch[28]~53 )) # (!Instr_ID_15 & ((!\pc_next_branch[28]~53 ) # (!nextPC_ID_29))))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [29]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[28]~53 ),
	.combout(\pc_next_branch[29]~54_combout ),
	.cout(\pc_next_branch[29]~55 ));
// synopsys translate_off
defparam \pc_next_branch[29]~54 .lut_mask = 16'h9617;
defparam \pc_next_branch[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \pc_next_branch[30]~56 (
// Equation(s):
// \pc_next_branch[30]~56_combout  = ((Instr_ID_15 $ (nextPC_ID_30 $ (!\pc_next_branch[29]~55 )))) # (GND)
// \pc_next_branch[30]~57  = CARRY((Instr_ID_15 & ((nextPC_ID_30) # (!\pc_next_branch[29]~55 ))) # (!Instr_ID_15 & (nextPC_ID_30 & !\pc_next_branch[29]~55 )))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [30]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[29]~55 ),
	.combout(\pc_next_branch[30]~56_combout ),
	.cout(\pc_next_branch[30]~57 ));
// synopsys translate_off
defparam \pc_next_branch[30]~56 .lut_mask = 16'h698E;
defparam \pc_next_branch[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N28
cycloneive_lcell_comb \pc_next_branch[31]~58 (
// Equation(s):
// \pc_next_branch[31]~58_combout  = nextPC_ID_31 $ (\pc_next_branch[30]~57  $ (Instr_ID_15))

	.dataa(gnd),
	.datab(\PR|nextPC_ID [31]),
	.datac(gnd),
	.datad(\PR|Instr_ID [15]),
	.cin(\pc_next_branch[30]~57 ),
	.combout(\pc_next_branch[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next_branch[31]~58 .lut_mask = 16'hC33C;
defparam \pc_next_branch[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \input_b~0 (
// Equation(s):
// \input_b~0_combout  = (!MemToReg_EX1 & (!Memwrite_ID1 & !Equal42))

	.dataa(MemToReg_EX),
	.datab(\PR|Memwrite_ID~q ),
	.datac(gnd),
	.datad(\HZ|Equal4~4_combout ),
	.cin(gnd),
	.combout(\input_b~0_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~0 .lut_mask = 16'h0011;
defparam \input_b~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \input_b~1 (
// Equation(s):
// \input_b~1_combout  = (\input_b~0_combout  & (!Equal4 & (!Equal41 & always0)))

	.dataa(\input_b~0_combout ),
	.datab(\HZ|Equal4~2_combout ),
	.datac(\HZ|Equal4~3_combout ),
	.datad(\HZ|always0~0_combout ),
	.cin(gnd),
	.combout(\input_b~1_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~1 .lut_mask = 16'h0200;
defparam \input_b~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \input_a~56 (
// Equation(s):
// \input_a~56_combout  = (MemToReg_MEM1 & ((ReadData_MEM_31))) # (!MemToReg_MEM1 & (CalcData_MEM_31))

	.dataa(\PR|CalcData_MEM [31]),
	.datab(\PR|ReadData_MEM [31]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~56_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~56 .lut_mask = 16'hCCAA;
defparam \input_a~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \output_RegWen_MEM~0 (
// Equation(s):
// \output_RegWen_MEM~0_combout  = (RegDst_MEM_0 & RegWen_MEM1)

	.dataa(gnd),
	.datab(gnd),
	.datac(\PR|RegDst_MEM [0]),
	.datad(\PR|RegWen_MEM~q ),
	.cin(gnd),
	.combout(\output_RegWen_MEM~0_combout ),
	.cout());
// synopsys translate_off
defparam \output_RegWen_MEM~0 .lut_mask = 16'hF000;
defparam \output_RegWen_MEM~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \output_RegWen_MEM~1 (
// Equation(s):
// \output_RegWen_MEM~1_combout  = (RegDst_MEM_4 & RegWen_MEM1)

	.dataa(\PR|RegDst_MEM [4]),
	.datab(\PR|RegWen_MEM~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\output_RegWen_MEM~1_combout ),
	.cout());
// synopsys translate_off
defparam \output_RegWen_MEM~1 .lut_mask = 16'h8888;
defparam \output_RegWen_MEM~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \input_b~2 (
// Equation(s):
// \input_b~2_combout  = (Memwrite_ID1) # ((!src2_hazard_t & !always01))

	.dataa(\HZ|src2_hazard_t~2_combout ),
	.datab(\PR|Memwrite_ID~q ),
	.datac(gnd),
	.datad(\HZ|always0~1_combout ),
	.cin(gnd),
	.combout(\input_b~2_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~2 .lut_mask = 16'hCCDD;
defparam \input_b~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \input_b~3 (
// Equation(s):
// \input_b~3_combout  = (!MemToReg_EX1) # (!MemToReg_MEM1)

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(MemToReg_EX),
	.cin(gnd),
	.combout(\input_b~3_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~3 .lut_mask = 16'h55FF;
defparam \input_b~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \input_b~4 (
// Equation(s):
// \input_b~4_combout  = (!Memwrite_ID1 & (!always01 & (\input_b~3_combout  & src2_hazard_t)))

	.dataa(\PR|Memwrite_ID~q ),
	.datab(\HZ|always0~1_combout ),
	.datac(\input_b~3_combout ),
	.datad(\HZ|src2_hazard_t~2_combout ),
	.cin(gnd),
	.combout(\input_b~4_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~4 .lut_mask = 16'h1000;
defparam \input_b~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \input_b~5 (
// Equation(s):
// \input_b~5_combout  = (ALUSrc2_ID_31 & ((\input_b~2_combout ) # ((\input_a~56_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_31 & (\input_a~56_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [31]),
	.datab(\input_a~56_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~5_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~5 .lut_mask = 16'hEAC0;
defparam \input_b~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \input_a~57 (
// Equation(s):
// \input_a~57_combout  = (!MemToReg_EX1 & (Instr_ID_23 $ (((!RegDst_EX_2) # (!RegWen_EX1)))))

	.dataa(\PR|RegWen_EX~q ),
	.datab(\PR|RegDst_EX [2]),
	.datac(\PR|Instr_ID [23]),
	.datad(MemToReg_EX),
	.cin(gnd),
	.combout(\input_a~57_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~57 .lut_mask = 16'h0087;
defparam \input_a~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \input_a~58 (
// Equation(s):
// \input_a~58_combout  = (!Equal01 & (\input_a~57_combout  & (!Equal0 & always02)))

	.dataa(\HZ|Equal0~3_combout ),
	.datab(\input_a~57_combout ),
	.datac(\HZ|Equal0~2_combout ),
	.datad(\HZ|always0~2_combout ),
	.cin(gnd),
	.combout(\input_a~58_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~58 .lut_mask = 16'h0400;
defparam \input_a~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \input_a~59 (
// Equation(s):
// \input_a~59_combout  = (\Equal22~0_combout  & (((Result_EX_31 & \input_a~58_combout )))) # (!\Equal22~0_combout  & ((ALUSrc1_ID_31) # ((Result_EX_31 & \input_a~58_combout ))))

	.dataa(\Equal22~0_combout ),
	.datab(\PR|ALUSrc1_ID [31]),
	.datac(Result_EX_31),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~59_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~59 .lut_mask = 16'hF444;
defparam \input_a~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \input_a~60 (
// Equation(s):
// \input_a~60_combout  = (always03 & (MemToReg_EX1)) # (!always03 & ((src1_hazard_t)))

	.dataa(MemToReg_EX),
	.datab(\HZ|always0~8_combout ),
	.datac(gnd),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\input_a~60_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~60 .lut_mask = 16'hBB88;
defparam \input_a~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \input_a~61 (
// Equation(s):
// \input_a~61_combout  = (\input_a~59_combout ) # ((\input_a~60_combout  & (\Equal24~0_combout  & \input_a~56_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~59_combout ),
	.datad(\input_a~56_combout ),
	.cin(gnd),
	.combout(\input_a~61_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~61 .lut_mask = 16'hF8F0;
defparam \input_a~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \input_b~6 (
// Equation(s):
// \input_b~6_combout  = (\input_b~5_combout ) # ((Result_EX_31 & \input_b~1_combout ))

	.dataa(Result_EX_31),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~5_combout ),
	.cin(gnd),
	.combout(\input_b~6_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~6 .lut_mask = 16'hFFA0;
defparam \input_b~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \input_a~62 (
// Equation(s):
// \input_a~62_combout  = (\Equal22~0_combout  & (Result_EX_30 & ((\input_a~58_combout )))) # (!\Equal22~0_combout  & ((ALUSrc1_ID_30) # ((Result_EX_30 & \input_a~58_combout ))))

	.dataa(\Equal22~0_combout ),
	.datab(Result_EX_30),
	.datac(\PR|ALUSrc1_ID [30]),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~62_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~62 .lut_mask = 16'hDC50;
defparam \input_a~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \input_b~7 (
// Equation(s):
// \input_b~7_combout  = (MemToReg_MEM1 & ((ReadData_MEM_30))) # (!MemToReg_MEM1 & (CalcData_MEM_30))

	.dataa(\PR|CalcData_MEM [30]),
	.datab(\PR|ReadData_MEM [30]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~7_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~7 .lut_mask = 16'hCCAA;
defparam \input_b~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \input_a~63 (
// Equation(s):
// \input_a~63_combout  = (\input_a~62_combout ) # ((\input_b~7_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_b~7_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~62_combout ),
	.datad(\input_a~60_combout ),
	.cin(gnd),
	.combout(\input_a~63_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~63 .lut_mask = 16'hF8F0;
defparam \input_a~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N24
cycloneive_lcell_comb \input_b~8 (
// Equation(s):
// \input_b~8_combout  = (\input_b~7_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_30 & \input_b~2_combout )))) # (!\input_b~7_combout  & (ALUSrc2_ID_30 & (\input_b~2_combout )))

	.dataa(\input_b~7_combout ),
	.datab(\PR|ALUSrc2_ID [30]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~8_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~8 .lut_mask = 16'hEAC0;
defparam \input_b~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N30
cycloneive_lcell_comb \input_b~9 (
// Equation(s):
// \input_b~9_combout  = (\input_b~8_combout ) # ((Result_EX_30 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_30),
	.datac(\input_b~1_combout ),
	.datad(\input_b~8_combout ),
	.cin(gnd),
	.combout(\input_b~9_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~9 .lut_mask = 16'hFFC0;
defparam \input_b~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \input_a~64 (
// Equation(s):
// \input_a~64_combout  = (ALUSrc1_ID_29 & (((Result_EX_29 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_29 & (Result_EX_29 & ((\input_a~58_combout ))))

	.dataa(\PR|ALUSrc1_ID [29]),
	.datab(Result_EX_29),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~64_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~64 .lut_mask = 16'hCE0A;
defparam \input_a~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \input_b~10 (
// Equation(s):
// \input_b~10_combout  = (MemToReg_MEM1 & (ReadData_MEM_29)) # (!MemToReg_MEM1 & ((CalcData_MEM_29)))

	.dataa(\PR|ReadData_MEM [29]),
	.datab(gnd),
	.datac(\PR|CalcData_MEM [29]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~10_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~10 .lut_mask = 16'hAAF0;
defparam \input_b~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \input_a~65 (
// Equation(s):
// \input_a~65_combout  = (\input_a~64_combout ) # ((\Equal24~0_combout  & (\input_b~10_combout  & \input_a~60_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_b~10_combout ),
	.datac(\input_a~64_combout ),
	.datad(\input_a~60_combout ),
	.cin(gnd),
	.combout(\input_a~65_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~65 .lut_mask = 16'hF8F0;
defparam \input_a~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N0
cycloneive_lcell_comb \input_b~11 (
// Equation(s):
// \input_b~11_combout  = (ALUSrc2_ID_29 & ((\input_b~2_combout ) # ((\input_b~10_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_29 & (\input_b~10_combout  & ((\input_b~4_combout ))))

	.dataa(\PR|ALUSrc2_ID [29]),
	.datab(\input_b~10_combout ),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~11_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~11 .lut_mask = 16'hECA0;
defparam \input_b~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N10
cycloneive_lcell_comb \input_b~12 (
// Equation(s):
// \input_b~12_combout  = (\input_b~11_combout ) # ((Result_EX_29 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_29),
	.datac(\input_b~1_combout ),
	.datad(\input_b~11_combout ),
	.cin(gnd),
	.combout(\input_b~12_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~12 .lut_mask = 16'hFFC0;
defparam \input_b~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \input_a~66 (
// Equation(s):
// \input_a~66_combout  = (ALUSrc1_ID_28 & (((Result_EX_28 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_28 & (Result_EX_28 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [28]),
	.datab(Result_EX_28),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~66_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~66 .lut_mask = 16'hC0EA;
defparam \input_a~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \input_b~13 (
// Equation(s):
// \input_b~13_combout  = (MemToReg_MEM1 & (ReadData_MEM_28)) # (!MemToReg_MEM1 & ((CalcData_MEM_28)))

	.dataa(\PR|ReadData_MEM [28]),
	.datab(gnd),
	.datac(\PR|CalcData_MEM [28]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~13_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~13 .lut_mask = 16'hAAF0;
defparam \input_b~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \input_a~67 (
// Equation(s):
// \input_a~67_combout  = (\input_a~66_combout ) # ((\Equal24~0_combout  & (\input_a~60_combout  & \input_b~13_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_a~60_combout ),
	.datac(\input_b~13_combout ),
	.datad(\input_a~66_combout ),
	.cin(gnd),
	.combout(\input_a~67_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~67 .lut_mask = 16'hFF80;
defparam \input_a~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \input_b~14 (
// Equation(s):
// \input_b~14_combout  = (ALUSrc2_ID_28 & ((\input_b~2_combout ) # ((\input_b~13_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_28 & (((\input_b~13_combout  & \input_b~4_combout ))))

	.dataa(\PR|ALUSrc2_ID [28]),
	.datab(\input_b~2_combout ),
	.datac(\input_b~13_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~14_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~14 .lut_mask = 16'hF888;
defparam \input_b~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N10
cycloneive_lcell_comb \input_b~15 (
// Equation(s):
// \input_b~15_combout  = (\input_b~14_combout ) # ((Result_EX_28 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_28),
	.datac(\input_b~1_combout ),
	.datad(\input_b~14_combout ),
	.cin(gnd),
	.combout(\input_b~15_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~15 .lut_mask = 16'hFFC0;
defparam \input_b~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \input_a~68 (
// Equation(s):
// \input_a~68_combout  = (\input_a~58_combout  & ((Result_EX_27) # ((ALUSrc1_ID_27 & !\Equal22~0_combout )))) # (!\input_a~58_combout  & (ALUSrc1_ID_27 & ((!\Equal22~0_combout ))))

	.dataa(\input_a~58_combout ),
	.datab(\PR|ALUSrc1_ID [27]),
	.datac(Result_EX_27),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~68_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~68 .lut_mask = 16'hA0EC;
defparam \input_a~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \input_b~16 (
// Equation(s):
// \input_b~16_combout  = (MemToReg_MEM1 & ((ReadData_MEM_27))) # (!MemToReg_MEM1 & (CalcData_MEM_27))

	.dataa(gnd),
	.datab(\PR|CalcData_MEM [27]),
	.datac(\PR|ReadData_MEM [27]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~16_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~16 .lut_mask = 16'hF0CC;
defparam \input_b~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \input_a~69 (
// Equation(s):
// \input_a~69_combout  = (\input_a~68_combout ) # ((\input_a~60_combout  & (\Equal24~0_combout  & \input_b~16_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_b~16_combout ),
	.datad(\input_a~68_combout ),
	.cin(gnd),
	.combout(\input_a~69_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~69 .lut_mask = 16'hFF80;
defparam \input_a~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \input_b~17 (
// Equation(s):
// \input_b~17_combout  = (\input_b~16_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_27 & \input_b~2_combout )))) # (!\input_b~16_combout  & (ALUSrc2_ID_27 & (\input_b~2_combout )))

	.dataa(\input_b~16_combout ),
	.datab(\PR|ALUSrc2_ID [27]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~17_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~17 .lut_mask = 16'hEAC0;
defparam \input_b~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \input_b~18 (
// Equation(s):
// \input_b~18_combout  = (\input_b~17_combout ) # ((Result_EX_27 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_27),
	.datac(\input_b~1_combout ),
	.datad(\input_b~17_combout ),
	.cin(gnd),
	.combout(\input_b~18_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~18 .lut_mask = 16'hFFC0;
defparam \input_b~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \input_a~70 (
// Equation(s):
// \input_a~70_combout  = (Result_EX_26 & ((\input_a~58_combout ) # ((ALUSrc1_ID_26 & !\Equal22~0_combout )))) # (!Result_EX_26 & (ALUSrc1_ID_26 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_26),
	.datab(\PR|ALUSrc1_ID [26]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~70_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~70 .lut_mask = 16'hA0EC;
defparam \input_a~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \input_b~19 (
// Equation(s):
// \input_b~19_combout  = (MemToReg_MEM1 & ((ReadData_MEM_26))) # (!MemToReg_MEM1 & (CalcData_MEM_26))

	.dataa(\PR|CalcData_MEM [26]),
	.datab(gnd),
	.datac(\PR|ReadData_MEM [26]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~19_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~19 .lut_mask = 16'hF0AA;
defparam \input_b~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \input_a~71 (
// Equation(s):
// \input_a~71_combout  = (\input_a~70_combout ) # ((\input_b~19_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_b~19_combout ),
	.datab(\input_a~70_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~60_combout ),
	.cin(gnd),
	.combout(\input_a~71_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~71 .lut_mask = 16'hECCC;
defparam \input_a~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \input_b~20 (
// Equation(s):
// \input_b~20_combout  = (\input_b~2_combout  & ((ALUSrc2_ID_26) # ((\input_b~19_combout  & \input_b~4_combout )))) # (!\input_b~2_combout  & (((\input_b~19_combout  & \input_b~4_combout ))))

	.dataa(\input_b~2_combout ),
	.datab(\PR|ALUSrc2_ID [26]),
	.datac(\input_b~19_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~20_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~20 .lut_mask = 16'hF888;
defparam \input_b~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \input_b~21 (
// Equation(s):
// \input_b~21_combout  = (\input_b~20_combout ) # ((Result_EX_26 & \input_b~1_combout ))

	.dataa(Result_EX_26),
	.datab(\input_b~1_combout ),
	.datac(\input_b~20_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\input_b~21_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~21 .lut_mask = 16'hF8F8;
defparam \input_b~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N4
cycloneive_lcell_comb \input_a~72 (
// Equation(s):
// \input_a~72_combout  = (ALUSrc1_ID_25 & (((Result_EX_25 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_25 & (Result_EX_25 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [25]),
	.datab(Result_EX_25),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~72_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~72 .lut_mask = 16'hC0EA;
defparam \input_a~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N18
cycloneive_lcell_comb \input_b~22 (
// Equation(s):
// \input_b~22_combout  = (MemToReg_MEM1 & (ReadData_MEM_25)) # (!MemToReg_MEM1 & ((CalcData_MEM_25)))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(gnd),
	.datac(\PR|ReadData_MEM [25]),
	.datad(\PR|CalcData_MEM [25]),
	.cin(gnd),
	.combout(\input_b~22_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~22 .lut_mask = 16'hF5A0;
defparam \input_b~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N0
cycloneive_lcell_comb \input_a~73 (
// Equation(s):
// \input_a~73_combout  = (\input_a~72_combout ) # ((\input_b~22_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_b~22_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~72_combout ),
	.datad(\input_a~60_combout ),
	.cin(gnd),
	.combout(\input_a~73_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~73 .lut_mask = 16'hF8F0;
defparam \input_a~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N2
cycloneive_lcell_comb \input_b~23 (
// Equation(s):
// \input_b~23_combout  = (ALUSrc2_ID_25 & ((\input_b~2_combout ) # ((\input_b~22_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_25 & (\input_b~22_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [25]),
	.datab(\input_b~22_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~23_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~23 .lut_mask = 16'hEAC0;
defparam \input_b~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N8
cycloneive_lcell_comb \input_b~24 (
// Equation(s):
// \input_b~24_combout  = (\input_b~23_combout ) # ((\input_b~1_combout  & Result_EX_25))

	.dataa(gnd),
	.datab(\input_b~1_combout ),
	.datac(Result_EX_25),
	.datad(\input_b~23_combout ),
	.cin(gnd),
	.combout(\input_b~24_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~24 .lut_mask = 16'hFFC0;
defparam \input_b~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N24
cycloneive_lcell_comb \input_a~74 (
// Equation(s):
// \input_a~74_combout  = (Result_EX_24 & ((\input_a~58_combout ) # ((ALUSrc1_ID_24 & !\Equal22~0_combout )))) # (!Result_EX_24 & (ALUSrc1_ID_24 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_24),
	.datab(\PR|ALUSrc1_ID [24]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~74_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~74 .lut_mask = 16'hA0EC;
defparam \input_a~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \input_b~25 (
// Equation(s):
// \input_b~25_combout  = (MemToReg_MEM1 & ((ReadData_MEM_24))) # (!MemToReg_MEM1 & (CalcData_MEM_24))

	.dataa(gnd),
	.datab(\PR|CalcData_MEM [24]),
	.datac(\PR|ReadData_MEM [24]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~25_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~25 .lut_mask = 16'hF0CC;
defparam \input_b~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N10
cycloneive_lcell_comb \input_a~75 (
// Equation(s):
// \input_a~75_combout  = (\input_a~74_combout ) # ((\Equal24~0_combout  & (\input_b~25_combout  & \input_a~60_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_b~25_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~74_combout ),
	.cin(gnd),
	.combout(\input_a~75_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~75 .lut_mask = 16'hFF80;
defparam \input_a~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N28
cycloneive_lcell_comb \input_b~26 (
// Equation(s):
// \input_b~26_combout  = (\input_b~25_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_24 & \input_b~2_combout )))) # (!\input_b~25_combout  & (ALUSrc2_ID_24 & (\input_b~2_combout )))

	.dataa(\input_b~25_combout ),
	.datab(\PR|ALUSrc2_ID [24]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~26_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~26 .lut_mask = 16'hEAC0;
defparam \input_b~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N6
cycloneive_lcell_comb \input_b~27 (
// Equation(s):
// \input_b~27_combout  = (\input_b~26_combout ) # ((\input_b~1_combout  & Result_EX_24))

	.dataa(\input_b~1_combout ),
	.datab(gnd),
	.datac(Result_EX_24),
	.datad(\input_b~26_combout ),
	.cin(gnd),
	.combout(\input_b~27_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~27 .lut_mask = 16'hFFA0;
defparam \input_b~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \input_a~76 (
// Equation(s):
// \input_a~76_combout  = (Result_EX_23 & ((\input_a~58_combout ) # ((ALUSrc1_ID_23 & !\Equal22~0_combout )))) # (!Result_EX_23 & (ALUSrc1_ID_23 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_23),
	.datab(\PR|ALUSrc1_ID [23]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~76_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~76 .lut_mask = 16'hA0EC;
defparam \input_a~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \input_b~28 (
// Equation(s):
// \input_b~28_combout  = (MemToReg_MEM1 & (ReadData_MEM_23)) # (!MemToReg_MEM1 & ((CalcData_MEM_23)))

	.dataa(\PR|ReadData_MEM [23]),
	.datab(\PR|CalcData_MEM [23]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\input_b~28_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~28 .lut_mask = 16'hACAC;
defparam \input_b~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \input_a~77 (
// Equation(s):
// \input_a~77_combout  = (\input_a~76_combout ) # ((\input_b~28_combout  & (\input_a~60_combout  & \Equal24~0_combout )))

	.dataa(\input_b~28_combout ),
	.datab(\input_a~60_combout ),
	.datac(\input_a~76_combout ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~77_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~77 .lut_mask = 16'hF8F0;
defparam \input_a~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \input_b~29 (
// Equation(s):
// \input_b~29_combout  = (\input_b~28_combout  & ((\input_b~4_combout ) # ((\input_b~2_combout  & ALUSrc2_ID_23)))) # (!\input_b~28_combout  & (\input_b~2_combout  & (ALUSrc2_ID_23)))

	.dataa(\input_b~28_combout ),
	.datab(\input_b~2_combout ),
	.datac(\PR|ALUSrc2_ID [23]),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~29_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~29 .lut_mask = 16'hEAC0;
defparam \input_b~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \input_b~30 (
// Equation(s):
// \input_b~30_combout  = (\input_b~29_combout ) # ((\input_b~1_combout  & Result_EX_23))

	.dataa(\input_b~1_combout ),
	.datab(Result_EX_23),
	.datac(gnd),
	.datad(\input_b~29_combout ),
	.cin(gnd),
	.combout(\input_b~30_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~30 .lut_mask = 16'hFF88;
defparam \input_b~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \input_a~78 (
// Equation(s):
// \input_a~78_combout  = (Result_EX_22 & ((\input_a~58_combout ) # ((ALUSrc1_ID_22 & !\Equal22~0_combout )))) # (!Result_EX_22 & (ALUSrc1_ID_22 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_22),
	.datab(\PR|ALUSrc1_ID [22]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~78_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~78 .lut_mask = 16'hA0EC;
defparam \input_a~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \input_b~31 (
// Equation(s):
// \input_b~31_combout  = (MemToReg_MEM1 & (ReadData_MEM_22)) # (!MemToReg_MEM1 & ((CalcData_MEM_22)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [22]),
	.datac(\PR|CalcData_MEM [22]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~31_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~31 .lut_mask = 16'hCCF0;
defparam \input_b~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \input_a~79 (
// Equation(s):
// \input_a~79_combout  = (\input_a~78_combout ) # ((\input_b~31_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_b~31_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~78_combout ),
	.cin(gnd),
	.combout(\input_a~79_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~79 .lut_mask = 16'hFF80;
defparam \input_a~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \input_b~32 (
// Equation(s):
// \input_b~32_combout  = (\input_b~31_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_22 & \input_b~2_combout )))) # (!\input_b~31_combout  & (ALUSrc2_ID_22 & ((\input_b~2_combout ))))

	.dataa(\input_b~31_combout ),
	.datab(\PR|ALUSrc2_ID [22]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~32_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~32 .lut_mask = 16'hECA0;
defparam \input_b~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \input_b~33 (
// Equation(s):
// \input_b~33_combout  = (\input_b~32_combout ) # ((Result_EX_22 & \input_b~1_combout ))

	.dataa(Result_EX_22),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~32_combout ),
	.cin(gnd),
	.combout(\input_b~33_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~33 .lut_mask = 16'hFFA0;
defparam \input_b~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \input_a~80 (
// Equation(s):
// \input_a~80_combout  = (Result_EX_21 & ((\input_a~58_combout ) # ((ALUSrc1_ID_21 & !\Equal22~0_combout )))) # (!Result_EX_21 & (ALUSrc1_ID_21 & (!\Equal22~0_combout )))

	.dataa(Result_EX_21),
	.datab(\PR|ALUSrc1_ID [21]),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~80_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~80 .lut_mask = 16'hAE0C;
defparam \input_a~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \input_b~34 (
// Equation(s):
// \input_b~34_combout  = (MemToReg_MEM1 & ((ReadData_MEM_21))) # (!MemToReg_MEM1 & (CalcData_MEM_21))

	.dataa(\PR|CalcData_MEM [21]),
	.datab(\PR|ReadData_MEM [21]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~34_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~34 .lut_mask = 16'hCCAA;
defparam \input_b~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \input_a~81 (
// Equation(s):
// \input_a~81_combout  = (\input_a~80_combout ) # ((\input_a~60_combout  & (\input_b~34_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_b~34_combout ),
	.datac(\input_a~80_combout ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~81_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~81 .lut_mask = 16'hF8F0;
defparam \input_a~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \input_b~35 (
// Equation(s):
// \input_b~35_combout  = (\input_b~34_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_21 & \input_b~2_combout )))) # (!\input_b~34_combout  & (ALUSrc2_ID_21 & (\input_b~2_combout )))

	.dataa(\input_b~34_combout ),
	.datab(\PR|ALUSrc2_ID [21]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~35_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~35 .lut_mask = 16'hEAC0;
defparam \input_b~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \input_b~36 (
// Equation(s):
// \input_b~36_combout  = (\input_b~35_combout ) # ((Result_EX_21 & \input_b~1_combout ))

	.dataa(Result_EX_21),
	.datab(\input_b~1_combout ),
	.datac(gnd),
	.datad(\input_b~35_combout ),
	.cin(gnd),
	.combout(\input_b~36_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~36 .lut_mask = 16'hFF88;
defparam \input_b~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \input_a~82 (
// Equation(s):
// \input_a~82_combout  = (ALUSrc1_ID_20 & (((Result_EX_20 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_20 & (Result_EX_20 & ((\input_a~58_combout ))))

	.dataa(\PR|ALUSrc1_ID [20]),
	.datab(Result_EX_20),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~82_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~82 .lut_mask = 16'hCE0A;
defparam \input_a~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \input_b~37 (
// Equation(s):
// \input_b~37_combout  = (MemToReg_MEM1 & ((ReadData_MEM_20))) # (!MemToReg_MEM1 & (CalcData_MEM_20))

	.dataa(\PR|CalcData_MEM [20]),
	.datab(\PR|ReadData_MEM [20]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~37_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~37 .lut_mask = 16'hCCAA;
defparam \input_b~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \input_a~83 (
// Equation(s):
// \input_a~83_combout  = (\input_a~82_combout ) # ((\input_a~60_combout  & (\input_b~37_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_b~37_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~82_combout ),
	.cin(gnd),
	.combout(\input_a~83_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~83 .lut_mask = 16'hFF80;
defparam \input_a~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \input_b~38 (
// Equation(s):
// \input_b~38_combout  = (ALUSrc2_ID_20 & ((\input_b~2_combout ) # ((\input_b~37_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_20 & (\input_b~37_combout  & ((\input_b~4_combout ))))

	.dataa(\PR|ALUSrc2_ID [20]),
	.datab(\input_b~37_combout ),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~38_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~38 .lut_mask = 16'hECA0;
defparam \input_b~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \input_b~39 (
// Equation(s):
// \input_b~39_combout  = (\input_b~38_combout ) # ((Result_EX_20 & \input_b~1_combout ))

	.dataa(Result_EX_20),
	.datab(\input_b~1_combout ),
	.datac(gnd),
	.datad(\input_b~38_combout ),
	.cin(gnd),
	.combout(\input_b~39_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~39 .lut_mask = 16'hFF88;
defparam \input_b~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \input_a~84 (
// Equation(s):
// \input_a~84_combout  = (Result_EX_19 & ((\input_a~58_combout ) # ((ALUSrc1_ID_19 & !\Equal22~0_combout )))) # (!Result_EX_19 & (ALUSrc1_ID_19 & (!\Equal22~0_combout )))

	.dataa(Result_EX_19),
	.datab(\PR|ALUSrc1_ID [19]),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~84_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~84 .lut_mask = 16'hAE0C;
defparam \input_a~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \input_b~40 (
// Equation(s):
// \input_b~40_combout  = (MemToReg_MEM1 & (ReadData_MEM_19)) # (!MemToReg_MEM1 & ((CalcData_MEM_19)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [19]),
	.datac(\PR|CalcData_MEM [19]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~40_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~40 .lut_mask = 16'hCCF0;
defparam \input_b~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \input_a~85 (
// Equation(s):
// \input_a~85_combout  = (\input_a~84_combout ) # ((\input_b~40_combout  & (\input_a~60_combout  & \Equal24~0_combout )))

	.dataa(\input_a~84_combout ),
	.datab(\input_b~40_combout ),
	.datac(\input_a~60_combout ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~85_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~85 .lut_mask = 16'hEAAA;
defparam \input_a~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \input_b~41 (
// Equation(s):
// \input_b~41_combout  = (ALUSrc2_ID_19 & ((\input_b~2_combout ) # ((\input_b~4_combout  & \input_b~40_combout )))) # (!ALUSrc2_ID_19 & (\input_b~4_combout  & (\input_b~40_combout )))

	.dataa(\PR|ALUSrc2_ID [19]),
	.datab(\input_b~4_combout ),
	.datac(\input_b~40_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~41_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~41 .lut_mask = 16'hEAC0;
defparam \input_b~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \input_b~42 (
// Equation(s):
// \input_b~42_combout  = (\input_b~41_combout ) # ((\input_b~1_combout  & Result_EX_19))

	.dataa(\input_b~1_combout ),
	.datab(Result_EX_19),
	.datac(gnd),
	.datad(\input_b~41_combout ),
	.cin(gnd),
	.combout(\input_b~42_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~42 .lut_mask = 16'hFF88;
defparam \input_b~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \input_a~86 (
// Equation(s):
// \input_a~86_combout  = (Result_EX_18 & ((\input_a~58_combout ) # ((ALUSrc1_ID_18 & !\Equal22~0_combout )))) # (!Result_EX_18 & (ALUSrc1_ID_18 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_18),
	.datab(\PR|ALUSrc1_ID [18]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~86_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~86 .lut_mask = 16'hA0EC;
defparam \input_a~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \input_b~43 (
// Equation(s):
// \input_b~43_combout  = (MemToReg_MEM1 & (ReadData_MEM_18)) # (!MemToReg_MEM1 & ((CalcData_MEM_18)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [18]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|CalcData_MEM [18]),
	.cin(gnd),
	.combout(\input_b~43_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~43 .lut_mask = 16'hCFC0;
defparam \input_b~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \input_a~87 (
// Equation(s):
// \input_a~87_combout  = (\input_a~86_combout ) # ((\input_b~43_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_a~86_combout ),
	.datab(\input_b~43_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~60_combout ),
	.cin(gnd),
	.combout(\input_a~87_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~87 .lut_mask = 16'hEAAA;
defparam \input_a~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \input_b~44 (
// Equation(s):
// \input_b~44_combout  = (\input_b~2_combout  & ((ALUSrc2_ID_18) # ((\input_b~43_combout  & \input_b~4_combout )))) # (!\input_b~2_combout  & (\input_b~43_combout  & ((\input_b~4_combout ))))

	.dataa(\input_b~2_combout ),
	.datab(\input_b~43_combout ),
	.datac(\PR|ALUSrc2_ID [18]),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~44_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~44 .lut_mask = 16'hECA0;
defparam \input_b~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \input_b~45 (
// Equation(s):
// \input_b~45_combout  = (\input_b~44_combout ) # ((Result_EX_18 & \input_b~1_combout ))

	.dataa(Result_EX_18),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~44_combout ),
	.cin(gnd),
	.combout(\input_b~45_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~45 .lut_mask = 16'hFFA0;
defparam \input_b~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \input_a~88 (
// Equation(s):
// \input_a~88_combout  = (Result_EX_17 & ((\input_a~58_combout ) # ((ALUSrc1_ID_17 & !\Equal22~0_combout )))) # (!Result_EX_17 & (ALUSrc1_ID_17 & (!\Equal22~0_combout )))

	.dataa(Result_EX_17),
	.datab(\PR|ALUSrc1_ID [17]),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~88_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~88 .lut_mask = 16'hAE0C;
defparam \input_a~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \input_b~46 (
// Equation(s):
// \input_b~46_combout  = (MemToReg_MEM1 & ((ReadData_MEM_17))) # (!MemToReg_MEM1 & (CalcData_MEM_17))

	.dataa(\PR|CalcData_MEM [17]),
	.datab(\PR|ReadData_MEM [17]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~46_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~46 .lut_mask = 16'hCCAA;
defparam \input_b~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \input_a~89 (
// Equation(s):
// \input_a~89_combout  = (\input_a~88_combout ) # ((\input_b~46_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_b~46_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~88_combout ),
	.cin(gnd),
	.combout(\input_a~89_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~89 .lut_mask = 16'hFF80;
defparam \input_a~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \input_b~47 (
// Equation(s):
// \input_b~47_combout  = (ALUSrc2_ID_17 & ((\input_b~2_combout ) # ((\input_b~46_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_17 & (\input_b~46_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [17]),
	.datab(\input_b~46_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~47_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~47 .lut_mask = 16'hEAC0;
defparam \input_b~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \input_b~48 (
// Equation(s):
// \input_b~48_combout  = (\input_b~47_combout ) # ((Result_EX_17 & \input_b~1_combout ))

	.dataa(Result_EX_17),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~47_combout ),
	.cin(gnd),
	.combout(\input_b~48_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~48 .lut_mask = 16'hFFA0;
defparam \input_b~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \input_a~90 (
// Equation(s):
// \input_a~90_combout  = (ALUSrc1_ID_16 & (((\input_a~58_combout  & Result_EX_16)) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_16 & (\input_a~58_combout  & (Result_EX_16)))

	.dataa(\PR|ALUSrc1_ID [16]),
	.datab(\input_a~58_combout ),
	.datac(Result_EX_16),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~90_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~90 .lut_mask = 16'hC0EA;
defparam \input_a~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \input_b~49 (
// Equation(s):
// \input_b~49_combout  = (MemToReg_MEM1 & (ReadData_MEM_16)) # (!MemToReg_MEM1 & ((CalcData_MEM_16)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [16]),
	.datac(\PR|CalcData_MEM [16]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~49_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~49 .lut_mask = 16'hCCF0;
defparam \input_b~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \input_a~91 (
// Equation(s):
// \input_a~91_combout  = (\input_a~90_combout ) # ((\input_a~60_combout  & (\Equal24~0_combout  & \input_b~49_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_b~49_combout ),
	.datad(\input_a~90_combout ),
	.cin(gnd),
	.combout(\input_a~91_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~91 .lut_mask = 16'hFF80;
defparam \input_a~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \input_b~50 (
// Equation(s):
// \input_b~50_combout  = (\input_b~49_combout  & ((\input_b~4_combout ) # ((\input_b~2_combout  & ALUSrc2_ID_16)))) # (!\input_b~49_combout  & (((\input_b~2_combout  & ALUSrc2_ID_16))))

	.dataa(\input_b~49_combout ),
	.datab(\input_b~4_combout ),
	.datac(\input_b~2_combout ),
	.datad(\PR|ALUSrc2_ID [16]),
	.cin(gnd),
	.combout(\input_b~50_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~50 .lut_mask = 16'hF888;
defparam \input_b~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \input_b~51 (
// Equation(s):
// \input_b~51_combout  = (\input_b~50_combout ) # ((Result_EX_16 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_16),
	.datac(\input_b~1_combout ),
	.datad(\input_b~50_combout ),
	.cin(gnd),
	.combout(\input_b~51_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~51 .lut_mask = 16'hFFC0;
defparam \input_b~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \input_a~92 (
// Equation(s):
// \input_a~92_combout  = (Result_EX_15 & ((\input_a~58_combout ) # ((ALUSrc1_ID_15 & !\Equal22~0_combout )))) # (!Result_EX_15 & (ALUSrc1_ID_15 & (!\Equal22~0_combout )))

	.dataa(Result_EX_15),
	.datab(\PR|ALUSrc1_ID [15]),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~92_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~92 .lut_mask = 16'hAE0C;
defparam \input_a~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \input_b~52 (
// Equation(s):
// \input_b~52_combout  = (MemToReg_MEM1 & ((ReadData_MEM_15))) # (!MemToReg_MEM1 & (CalcData_MEM_15))

	.dataa(\PR|CalcData_MEM [15]),
	.datab(gnd),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|ReadData_MEM [15]),
	.cin(gnd),
	.combout(\input_b~52_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~52 .lut_mask = 16'hFA0A;
defparam \input_b~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N20
cycloneive_lcell_comb \input_a~93 (
// Equation(s):
// \input_a~93_combout  = (\input_a~92_combout ) # ((\input_a~60_combout  & (\input_b~52_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_b~52_combout ),
	.datac(\input_a~92_combout ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~93_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~93 .lut_mask = 16'hF8F0;
defparam \input_a~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \input_b~53 (
// Equation(s):
// \input_b~53_combout  = (ALUSrc2_ID_15 & ((\input_b~2_combout ) # ((\input_b~52_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_15 & (\input_b~52_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [15]),
	.datab(\input_b~52_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~53_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~53 .lut_mask = 16'hEAC0;
defparam \input_b~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N22
cycloneive_lcell_comb \input_b~54 (
// Equation(s):
// \input_b~54_combout  = (\input_b~53_combout ) # ((\input_b~1_combout  & Result_EX_15))

	.dataa(\input_b~1_combout ),
	.datab(gnd),
	.datac(Result_EX_15),
	.datad(\input_b~53_combout ),
	.cin(gnd),
	.combout(\input_b~54_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~54 .lut_mask = 16'hFFA0;
defparam \input_b~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N12
cycloneive_lcell_comb \input_a~94 (
// Equation(s):
// \input_a~94_combout  = (ALUSrc1_ID_14 & (((Result_EX_14 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_14 & (Result_EX_14 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [14]),
	.datab(Result_EX_14),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~94_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~94 .lut_mask = 16'hC0EA;
defparam \input_a~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N26
cycloneive_lcell_comb \input_b~55 (
// Equation(s):
// \input_b~55_combout  = (MemToReg_MEM1 & ((ReadData_MEM_14))) # (!MemToReg_MEM1 & (CalcData_MEM_14))

	.dataa(\PR|CalcData_MEM [14]),
	.datab(gnd),
	.datac(\PR|ReadData_MEM [14]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_b~55_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~55 .lut_mask = 16'hF0AA;
defparam \input_b~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N6
cycloneive_lcell_comb \input_a~95 (
// Equation(s):
// \input_a~95_combout  = (\input_a~94_combout ) # ((\input_b~55_combout  & (\input_a~60_combout  & \Equal24~0_combout )))

	.dataa(\input_b~55_combout ),
	.datab(\input_a~60_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~94_combout ),
	.cin(gnd),
	.combout(\input_a~95_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~95 .lut_mask = 16'hFF80;
defparam \input_a~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N10
cycloneive_lcell_comb \input_b~56 (
// Equation(s):
// \input_b~56_combout  = (\input_b~55_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_14 & \input_b~2_combout )))) # (!\input_b~55_combout  & (ALUSrc2_ID_14 & ((\input_b~2_combout ))))

	.dataa(\input_b~55_combout ),
	.datab(\PR|ALUSrc2_ID [14]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~56_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~56 .lut_mask = 16'hECA0;
defparam \input_b~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N8
cycloneive_lcell_comb \input_b~57 (
// Equation(s):
// \input_b~57_combout  = (\input_b~56_combout ) # ((\input_b~1_combout  & Result_EX_14))

	.dataa(\input_b~1_combout ),
	.datab(Result_EX_14),
	.datac(gnd),
	.datad(\input_b~56_combout ),
	.cin(gnd),
	.combout(\input_b~57_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~57 .lut_mask = 16'hFF88;
defparam \input_b~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N20
cycloneive_lcell_comb \input_a~96 (
// Equation(s):
// \input_a~96_combout  = (MemToReg_MEM1 & ((ReadData_MEM_13))) # (!MemToReg_MEM1 & (CalcData_MEM_13))

	.dataa(\PR|CalcData_MEM [13]),
	.datab(gnd),
	.datac(\PR|ReadData_MEM [13]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~96_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~96 .lut_mask = 16'hF0AA;
defparam \input_a~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N18
cycloneive_lcell_comb \input_b~58 (
// Equation(s):
// \input_b~58_combout  = (\input_a~96_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_13 & \input_b~2_combout )))) # (!\input_a~96_combout  & (ALUSrc2_ID_13 & ((\input_b~2_combout ))))

	.dataa(\input_a~96_combout ),
	.datab(\PR|ALUSrc2_ID [13]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~58_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~58 .lut_mask = 16'hECA0;
defparam \input_b~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N20
cycloneive_lcell_comb \input_b~59 (
// Equation(s):
// \input_b~59_combout  = (\input_b~58_combout ) # ((Result_EX_13 & \input_b~1_combout ))

	.dataa(Result_EX_13),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~58_combout ),
	.cin(gnd),
	.combout(\input_b~59_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~59 .lut_mask = 16'hFFA0;
defparam \input_b~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N26
cycloneive_lcell_comb \input_a~97 (
// Equation(s):
// \input_a~97_combout  = (ALUSrc1_ID_13 & (((Result_EX_13 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_13 & (Result_EX_13 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [13]),
	.datab(Result_EX_13),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~97_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~97 .lut_mask = 16'hC0EA;
defparam \input_a~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \input_a~98 (
// Equation(s):
// \input_a~98_combout  = (\input_a~97_combout ) # ((\input_a~60_combout  & (\input_a~96_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_a~96_combout ),
	.datac(\input_a~97_combout ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~98_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~98 .lut_mask = 16'hF8F0;
defparam \input_a~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N12
cycloneive_lcell_comb \input_a~99 (
// Equation(s):
// \input_a~99_combout  = (MemToReg_MEM1 & (ReadData_MEM_12)) # (!MemToReg_MEM1 & ((CalcData_MEM_12)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [12]),
	.datac(\PR|CalcData_MEM [12]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~99_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~99 .lut_mask = 16'hCCF0;
defparam \input_a~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N18
cycloneive_lcell_comb \input_b~60 (
// Equation(s):
// \input_b~60_combout  = (\input_a~99_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_12 & \input_b~2_combout )))) # (!\input_a~99_combout  & (ALUSrc2_ID_12 & (\input_b~2_combout )))

	.dataa(\input_a~99_combout ),
	.datab(\PR|ALUSrc2_ID [12]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~60_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~60 .lut_mask = 16'hEAC0;
defparam \input_b~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N0
cycloneive_lcell_comb \input_b~61 (
// Equation(s):
// \input_b~61_combout  = (\input_b~60_combout ) # ((Result_EX_12 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_12),
	.datac(\input_b~1_combout ),
	.datad(\input_b~60_combout ),
	.cin(gnd),
	.combout(\input_b~61_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~61 .lut_mask = 16'hFFC0;
defparam \input_b~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N14
cycloneive_lcell_comb \input_a~100 (
// Equation(s):
// \input_a~100_combout  = (ALUSrc1_ID_12 & (((Result_EX_12 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_12 & (Result_EX_12 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [12]),
	.datab(Result_EX_12),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~100_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~100 .lut_mask = 16'hC0EA;
defparam \input_a~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N20
cycloneive_lcell_comb \input_a~101 (
// Equation(s):
// \input_a~101_combout  = (\input_a~100_combout ) # ((\Equal24~0_combout  & (\input_a~60_combout  & \input_a~99_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_a~100_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~99_combout ),
	.cin(gnd),
	.combout(\input_a~101_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~101 .lut_mask = 16'hECCC;
defparam \input_a~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N26
cycloneive_lcell_comb \input_a~102 (
// Equation(s):
// \input_a~102_combout  = (MemToReg_MEM1 & (ReadData_MEM_11)) # (!MemToReg_MEM1 & ((CalcData_MEM_11)))

	.dataa(\PR|ReadData_MEM [11]),
	.datab(gnd),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|CalcData_MEM [11]),
	.cin(gnd),
	.combout(\input_a~102_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~102 .lut_mask = 16'hAFA0;
defparam \input_a~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N12
cycloneive_lcell_comb \input_b~62 (
// Equation(s):
// \input_b~62_combout  = (ALUSrc2_ID_11 & ((\input_b~2_combout ) # ((\input_a~102_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_11 & (\input_a~102_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [11]),
	.datab(\input_a~102_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~62_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~62 .lut_mask = 16'hEAC0;
defparam \input_b~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N14
cycloneive_lcell_comb \input_b~63 (
// Equation(s):
// \input_b~63_combout  = (\input_b~62_combout ) # ((\input_b~1_combout  & Result_EX_11))

	.dataa(\input_b~1_combout ),
	.datab(gnd),
	.datac(Result_EX_11),
	.datad(\input_b~62_combout ),
	.cin(gnd),
	.combout(\input_b~63_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~63 .lut_mask = 16'hFFA0;
defparam \input_b~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N12
cycloneive_lcell_comb \input_a~103 (
// Equation(s):
// \input_a~103_combout  = (Result_EX_11 & ((\input_a~58_combout ) # ((ALUSrc1_ID_11 & !\Equal22~0_combout )))) # (!Result_EX_11 & (ALUSrc1_ID_11 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_11),
	.datab(\PR|ALUSrc1_ID [11]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~103_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~103 .lut_mask = 16'hA0EC;
defparam \input_a~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N10
cycloneive_lcell_comb \input_a~104 (
// Equation(s):
// \input_a~104_combout  = (\input_a~103_combout ) # ((\input_a~102_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_a~102_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~103_combout ),
	.cin(gnd),
	.combout(\input_a~104_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~104 .lut_mask = 16'hFF80;
defparam \input_a~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N0
cycloneive_lcell_comb \input_a~105 (
// Equation(s):
// \input_a~105_combout  = (MemToReg_MEM1 & ((ReadData_MEM_10))) # (!MemToReg_MEM1 & (CalcData_MEM_10))

	.dataa(gnd),
	.datab(\PR|CalcData_MEM [10]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|ReadData_MEM [10]),
	.cin(gnd),
	.combout(\input_a~105_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~105 .lut_mask = 16'hFC0C;
defparam \input_a~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N6
cycloneive_lcell_comb \input_b~64 (
// Equation(s):
// \input_b~64_combout  = (\input_a~105_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_10 & \input_b~2_combout )))) # (!\input_a~105_combout  & (ALUSrc2_ID_10 & ((\input_b~2_combout ))))

	.dataa(\input_a~105_combout ),
	.datab(\PR|ALUSrc2_ID [10]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~64_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~64 .lut_mask = 16'hECA0;
defparam \input_b~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N4
cycloneive_lcell_comb \input_b~65 (
// Equation(s):
// \input_b~65_combout  = (\input_b~64_combout ) # ((\input_b~1_combout  & Result_EX_10))

	.dataa(\input_b~1_combout ),
	.datab(gnd),
	.datac(Result_EX_10),
	.datad(\input_b~64_combout ),
	.cin(gnd),
	.combout(\input_b~65_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~65 .lut_mask = 16'hFFA0;
defparam \input_b~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N18
cycloneive_lcell_comb \input_a~106 (
// Equation(s):
// \input_a~106_combout  = (ALUSrc1_ID_10 & (((Result_EX_10 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_10 & (Result_EX_10 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [10]),
	.datab(Result_EX_10),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~106_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~106 .lut_mask = 16'hC0EA;
defparam \input_a~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N16
cycloneive_lcell_comb \input_a~107 (
// Equation(s):
// \input_a~107_combout  = (\input_a~106_combout ) # ((\input_a~105_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_a~105_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~106_combout ),
	.cin(gnd),
	.combout(\input_a~107_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~107 .lut_mask = 16'hFF80;
defparam \input_a~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \input_a~108 (
// Equation(s):
// \input_a~108_combout  = (MemToReg_MEM1 & (ReadData_MEM_9)) # (!MemToReg_MEM1 & ((CalcData_MEM_9)))

	.dataa(\PR|ReadData_MEM [9]),
	.datab(gnd),
	.datac(\PR|CalcData_MEM [9]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~108_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~108 .lut_mask = 16'hAAF0;
defparam \input_a~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N16
cycloneive_lcell_comb \input_b~66 (
// Equation(s):
// \input_b~66_combout  = (\input_a~108_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_9 & \input_b~2_combout )))) # (!\input_a~108_combout  & (ALUSrc2_ID_9 & ((\input_b~2_combout ))))

	.dataa(\input_a~108_combout ),
	.datab(\PR|ALUSrc2_ID [9]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~66_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~66 .lut_mask = 16'hECA0;
defparam \input_b~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N2
cycloneive_lcell_comb \input_b~67 (
// Equation(s):
// \input_b~67_combout  = (\input_b~66_combout ) # ((Result_EX_9 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_9),
	.datac(\input_b~1_combout ),
	.datad(\input_b~66_combout ),
	.cin(gnd),
	.combout(\input_b~67_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~67 .lut_mask = 16'hFFC0;
defparam \input_b~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N12
cycloneive_lcell_comb \input_a~109 (
// Equation(s):
// \input_a~109_combout  = (ALUSrc1_ID_9 & (((Result_EX_9 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_9 & (Result_EX_9 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [9]),
	.datab(Result_EX_9),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~109_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~109 .lut_mask = 16'hC0EA;
defparam \input_a~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N30
cycloneive_lcell_comb \input_a~110 (
// Equation(s):
// \input_a~110_combout  = (\input_a~109_combout ) # ((\input_a~108_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_a~108_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~109_combout ),
	.cin(gnd),
	.combout(\input_a~110_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~110 .lut_mask = 16'hFF80;
defparam \input_a~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \input_a~111 (
// Equation(s):
// \input_a~111_combout  = (MemToReg_MEM1 & (ReadData_MEM_8)) # (!MemToReg_MEM1 & ((CalcData_MEM_8)))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|ReadData_MEM [8]),
	.datac(gnd),
	.datad(\PR|CalcData_MEM [8]),
	.cin(gnd),
	.combout(\input_a~111_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~111 .lut_mask = 16'hDD88;
defparam \input_a~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N10
cycloneive_lcell_comb \input_b~68 (
// Equation(s):
// \input_b~68_combout  = (ALUSrc2_ID_8 & ((\input_b~2_combout ) # ((\input_a~111_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_8 & (\input_a~111_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [8]),
	.datab(\input_a~111_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~68_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~68 .lut_mask = 16'hEAC0;
defparam \input_b~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \input_b~69 (
// Equation(s):
// \input_b~69_combout  = (\input_b~68_combout ) # ((\input_b~1_combout  & Result_EX_8))

	.dataa(\input_b~1_combout ),
	.datab(Result_EX_8),
	.datac(gnd),
	.datad(\input_b~68_combout ),
	.cin(gnd),
	.combout(\input_b~69_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~69 .lut_mask = 16'hFF88;
defparam \input_b~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \input_a~112 (
// Equation(s):
// \input_a~112_combout  = (Result_EX_8 & ((\input_a~58_combout ) # ((ALUSrc1_ID_8 & !\Equal22~0_combout )))) # (!Result_EX_8 & (ALUSrc1_ID_8 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_8),
	.datab(\PR|ALUSrc1_ID [8]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~112_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~112 .lut_mask = 16'hA0EC;
defparam \input_a~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \input_a~113 (
// Equation(s):
// \input_a~113_combout  = (\input_a~112_combout ) # ((\input_a~111_combout  & (\input_a~60_combout  & \Equal24~0_combout )))

	.dataa(\input_a~111_combout ),
	.datab(\input_a~60_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~112_combout ),
	.cin(gnd),
	.combout(\input_a~113_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~113 .lut_mask = 16'hFF80;
defparam \input_a~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \input_a~114 (
// Equation(s):
// \input_a~114_combout  = (MemToReg_MEM1 & (ReadData_MEM_7)) # (!MemToReg_MEM1 & ((CalcData_MEM_7)))

	.dataa(\PR|ReadData_MEM [7]),
	.datab(\PR|CalcData_MEM [7]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~114_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~114 .lut_mask = 16'hAACC;
defparam \input_a~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \input_b~70 (
// Equation(s):
// \input_b~70_combout  = (\input_a~114_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_7 & \input_b~2_combout )))) # (!\input_a~114_combout  & (ALUSrc2_ID_7 & (\input_b~2_combout )))

	.dataa(\input_a~114_combout ),
	.datab(\PR|ALUSrc2_ID [7]),
	.datac(\input_b~2_combout ),
	.datad(\input_b~4_combout ),
	.cin(gnd),
	.combout(\input_b~70_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~70 .lut_mask = 16'hEAC0;
defparam \input_b~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \input_b~71 (
// Equation(s):
// \input_b~71_combout  = (\input_b~70_combout ) # ((Result_EX_7 & \input_b~1_combout ))

	.dataa(Result_EX_7),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(\input_b~70_combout ),
	.cin(gnd),
	.combout(\input_b~71_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~71 .lut_mask = 16'hFFA0;
defparam \input_b~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \input_a~115 (
// Equation(s):
// \input_a~115_combout  = (Result_EX_7 & ((\input_a~58_combout ) # ((ALUSrc1_ID_7 & !\Equal22~0_combout )))) # (!Result_EX_7 & (ALUSrc1_ID_7 & ((!\Equal22~0_combout ))))

	.dataa(Result_EX_7),
	.datab(\PR|ALUSrc1_ID [7]),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~115_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~115 .lut_mask = 16'hA0EC;
defparam \input_a~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \input_a~116 (
// Equation(s):
// \input_a~116_combout  = (\input_a~115_combout ) # ((\input_a~114_combout  & (\Equal24~0_combout  & \input_a~60_combout )))

	.dataa(\input_a~114_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~115_combout ),
	.cin(gnd),
	.combout(\input_a~116_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~116 .lut_mask = 16'hFF80;
defparam \input_a~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \input_a~117 (
// Equation(s):
// \input_a~117_combout  = (MemToReg_MEM1 & ((ReadData_MEM_6))) # (!MemToReg_MEM1 & (CalcData_MEM_6))

	.dataa(\PR|CalcData_MEM [6]),
	.datab(gnd),
	.datac(\PR|ReadData_MEM [6]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~117_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~117 .lut_mask = 16'hF0AA;
defparam \input_a~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \input_b~72 (
// Equation(s):
// \input_b~72_combout  = (\input_a~117_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_6 & \input_b~2_combout )))) # (!\input_a~117_combout  & (ALUSrc2_ID_6 & ((\input_b~2_combout ))))

	.dataa(\input_a~117_combout ),
	.datab(\PR|ALUSrc2_ID [6]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~72_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~72 .lut_mask = 16'hECA0;
defparam \input_b~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \input_b~73 (
// Equation(s):
// \input_b~73_combout  = (\input_b~72_combout ) # ((Result_EX_6 & \input_b~1_combout ))

	.dataa(Result_EX_6),
	.datab(\input_b~1_combout ),
	.datac(gnd),
	.datad(\input_b~72_combout ),
	.cin(gnd),
	.combout(\input_b~73_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~73 .lut_mask = 16'hFF88;
defparam \input_b~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N12
cycloneive_lcell_comb \input_a~118 (
// Equation(s):
// \input_a~118_combout  = (Result_EX_6 & ((\input_a~58_combout ) # ((ALUSrc1_ID_6 & !\Equal22~0_combout )))) # (!Result_EX_6 & (ALUSrc1_ID_6 & (!\Equal22~0_combout )))

	.dataa(Result_EX_6),
	.datab(\PR|ALUSrc1_ID [6]),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~118_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~118 .lut_mask = 16'hAE0C;
defparam \input_a~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N30
cycloneive_lcell_comb \input_a~119 (
// Equation(s):
// \input_a~119_combout  = (\input_a~118_combout ) # ((\input_a~60_combout  & (\input_a~117_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_a~117_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~118_combout ),
	.cin(gnd),
	.combout(\input_a~119_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~119 .lut_mask = 16'hFF80;
defparam \input_a~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \input_a~120 (
// Equation(s):
// \input_a~120_combout  = (MemToReg_MEM1 & (ReadData_MEM_5)) # (!MemToReg_MEM1 & ((CalcData_MEM_5)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [5]),
	.datac(\PR|CalcData_MEM [5]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~120_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~120 .lut_mask = 16'hCCF0;
defparam \input_a~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \input_b~74 (
// Equation(s):
// \input_b~74_combout  = (\input_a~120_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_5 & \input_b~2_combout )))) # (!\input_a~120_combout  & (ALUSrc2_ID_5 & ((\input_b~2_combout ))))

	.dataa(\input_a~120_combout ),
	.datab(\PR|ALUSrc2_ID [5]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~74_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~74 .lut_mask = 16'hECA0;
defparam \input_b~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \input_b~75 (
// Equation(s):
// \input_b~75_combout  = (\input_b~74_combout ) # ((Result_EX_5 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_5),
	.datac(\input_b~1_combout ),
	.datad(\input_b~74_combout ),
	.cin(gnd),
	.combout(\input_b~75_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~75 .lut_mask = 16'hFFC0;
defparam \input_b~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \input_a~121 (
// Equation(s):
// \input_a~121_combout  = (ALUSrc1_ID_5 & (((Result_EX_5 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_5 & (Result_EX_5 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [5]),
	.datab(Result_EX_5),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~121_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~121 .lut_mask = 16'hC0EA;
defparam \input_a~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \input_a~122 (
// Equation(s):
// \input_a~122_combout  = (\input_a~121_combout ) # ((\input_a~120_combout  & (\input_a~60_combout  & \Equal24~0_combout )))

	.dataa(\input_a~120_combout ),
	.datab(\input_a~60_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~121_combout ),
	.cin(gnd),
	.combout(\input_a~122_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~122 .lut_mask = 16'hFF80;
defparam \input_a~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N16
cycloneive_lcell_comb \input_a~123 (
// Equation(s):
// \input_a~123_combout  = (MemToReg_MEM1 & ((ReadData_MEM_4))) # (!MemToReg_MEM1 & (CalcData_MEM_4))

	.dataa(\PR|CalcData_MEM [4]),
	.datab(\PR|ReadData_MEM [4]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~123_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~123 .lut_mask = 16'hCCAA;
defparam \input_a~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N28
cycloneive_lcell_comb \input_b~76 (
// Equation(s):
// \input_b~76_combout  = (\input_a~123_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_4 & \input_b~2_combout )))) # (!\input_a~123_combout  & (ALUSrc2_ID_4 & ((\input_b~2_combout ))))

	.dataa(\input_a~123_combout ),
	.datab(\PR|ALUSrc2_ID [4]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~76_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~76 .lut_mask = 16'hECA0;
defparam \input_b~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N10
cycloneive_lcell_comb \input_b~77 (
// Equation(s):
// \input_b~77_combout  = (\input_b~76_combout ) # ((\input_b~1_combout  & Result_EX_4))

	.dataa(\input_b~1_combout ),
	.datab(gnd),
	.datac(Result_EX_4),
	.datad(\input_b~76_combout ),
	.cin(gnd),
	.combout(\input_b~77_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~77 .lut_mask = 16'hFFA0;
defparam \input_b~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N10
cycloneive_lcell_comb \input_a~124 (
// Equation(s):
// \input_a~124_combout  = (ALUSrc1_ID_4 & (((Result_EX_4 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_4 & (Result_EX_4 & ((\input_a~58_combout ))))

	.dataa(\PR|ALUSrc1_ID [4]),
	.datab(Result_EX_4),
	.datac(\Equal22~0_combout ),
	.datad(\input_a~58_combout ),
	.cin(gnd),
	.combout(\input_a~124_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~124 .lut_mask = 16'hCE0A;
defparam \input_a~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N20
cycloneive_lcell_comb \input_a~125 (
// Equation(s):
// \input_a~125_combout  = (\input_a~124_combout ) # ((\input_a~60_combout  & (\input_a~123_combout  & \Equal24~0_combout )))

	.dataa(\input_a~60_combout ),
	.datab(\input_a~123_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\input_a~124_combout ),
	.cin(gnd),
	.combout(\input_a~125_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~125 .lut_mask = 16'hFF80;
defparam \input_a~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \input_a~126 (
// Equation(s):
// \input_a~126_combout  = (MemToReg_MEM1 & (ReadData_MEM_3)) # (!MemToReg_MEM1 & ((CalcData_MEM_3)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [3]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|CalcData_MEM [3]),
	.cin(gnd),
	.combout(\input_a~126_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~126 .lut_mask = 16'hCFC0;
defparam \input_a~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \input_b~78 (
// Equation(s):
// \input_b~78_combout  = (\input_a~126_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_3 & \input_b~2_combout )))) # (!\input_a~126_combout  & (ALUSrc2_ID_3 & ((\input_b~2_combout ))))

	.dataa(\input_a~126_combout ),
	.datab(\PR|ALUSrc2_ID [3]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~78_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~78 .lut_mask = 16'hECA0;
defparam \input_b~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \input_b~79 (
// Equation(s):
// \input_b~79_combout  = (\input_b~78_combout ) # ((Result_EX_3 & \input_b~1_combout ))

	.dataa(Result_EX_3),
	.datab(\input_b~1_combout ),
	.datac(gnd),
	.datad(\input_b~78_combout ),
	.cin(gnd),
	.combout(\input_b~79_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~79 .lut_mask = 16'hFF88;
defparam \input_b~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N18
cycloneive_lcell_comb \input_a~127 (
// Equation(s):
// \input_a~127_combout  = (ALUSrc1_ID_3 & (((Result_EX_3 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_3 & (Result_EX_3 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [3]),
	.datab(Result_EX_3),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~127_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~127 .lut_mask = 16'hC0EA;
defparam \input_a~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N16
cycloneive_lcell_comb \input_a~128 (
// Equation(s):
// \input_a~128_combout  = (\input_a~127_combout ) # ((\Equal24~0_combout  & (\input_a~126_combout  & \input_a~60_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_a~126_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~127_combout ),
	.cin(gnd),
	.combout(\input_a~128_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~128 .lut_mask = 16'hFF80;
defparam \input_a~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N8
cycloneive_lcell_comb \input_a~129 (
// Equation(s):
// \input_a~129_combout  = (MemToReg_MEM1 & ((ReadData_MEM_2))) # (!MemToReg_MEM1 & (CalcData_MEM_2))

	.dataa(\PR|CalcData_MEM [2]),
	.datab(gnd),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|ReadData_MEM [2]),
	.cin(gnd),
	.combout(\input_a~129_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~129 .lut_mask = 16'hFA0A;
defparam \input_a~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N6
cycloneive_lcell_comb \input_b~80 (
// Equation(s):
// \input_b~80_combout  = (ALUSrc2_ID_2 & ((\input_b~2_combout ) # ((\input_a~129_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_2 & (\input_a~129_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [2]),
	.datab(\input_a~129_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~80_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~80 .lut_mask = 16'hEAC0;
defparam \input_b~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N20
cycloneive_lcell_comb \input_b~81 (
// Equation(s):
// \input_b~81_combout  = (\input_b~80_combout ) # ((\input_b~1_combout  & Result_EX_2))

	.dataa(\input_b~1_combout ),
	.datab(Result_EX_2),
	.datac(gnd),
	.datad(\input_b~80_combout ),
	.cin(gnd),
	.combout(\input_b~81_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~81 .lut_mask = 16'hFF88;
defparam \input_b~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N2
cycloneive_lcell_comb \input_a~130 (
// Equation(s):
// \input_a~130_combout  = (ALUSrc1_ID_2 & (((Result_EX_2 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_2 & (Result_EX_2 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [2]),
	.datab(Result_EX_2),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~130_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~130 .lut_mask = 16'hC0EA;
defparam \input_a~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \input_a~131 (
// Equation(s):
// \input_a~131_combout  = (\input_a~130_combout ) # ((\Equal24~0_combout  & (\input_a~129_combout  & \input_a~60_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_a~129_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~130_combout ),
	.cin(gnd),
	.combout(\input_a~131_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~131 .lut_mask = 16'hFF80;
defparam \input_a~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \input_b~82 (
// Equation(s):
// \input_b~82_combout  = (ALUSrc2_ID_1 & ((\input_b~2_combout ) # ((\input_a~132_combout  & \input_b~4_combout )))) # (!ALUSrc2_ID_1 & (\input_a~132_combout  & (\input_b~4_combout )))

	.dataa(\PR|ALUSrc2_ID [1]),
	.datab(\input_a~132_combout ),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~82_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~82 .lut_mask = 16'hEAC0;
defparam \input_b~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N30
cycloneive_lcell_comb \input_b~83 (
// Equation(s):
// \input_b~83_combout  = (\input_b~82_combout ) # ((Result_EX_1 & \input_b~1_combout ))

	.dataa(gnd),
	.datab(Result_EX_1),
	.datac(\input_b~82_combout ),
	.datad(\input_b~1_combout ),
	.cin(gnd),
	.combout(\input_b~83_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~83 .lut_mask = 16'hFCF0;
defparam \input_b~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N0
cycloneive_lcell_comb \input_a~133 (
// Equation(s):
// \input_a~133_combout  = (ALUSrc1_ID_1 & (((Result_EX_1 & \input_a~58_combout )) # (!\Equal22~0_combout ))) # (!ALUSrc1_ID_1 & (Result_EX_1 & (\input_a~58_combout )))

	.dataa(\PR|ALUSrc1_ID [1]),
	.datab(Result_EX_1),
	.datac(\input_a~58_combout ),
	.datad(\Equal22~0_combout ),
	.cin(gnd),
	.combout(\input_a~133_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~133 .lut_mask = 16'hC0EA;
defparam \input_a~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N26
cycloneive_lcell_comb \input_a~134 (
// Equation(s):
// \input_a~134_combout  = (\input_a~133_combout ) # ((\Equal24~0_combout  & (\input_a~132_combout  & \input_a~60_combout )))

	.dataa(\Equal24~0_combout ),
	.datab(\input_a~132_combout ),
	.datac(\input_a~60_combout ),
	.datad(\input_a~133_combout ),
	.cin(gnd),
	.combout(\input_a~134_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~134 .lut_mask = 16'hFF80;
defparam \input_a~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \input_b~84 (
// Equation(s):
// \input_b~84_combout  = (\input_a~135_combout  & ((\input_b~4_combout ) # ((ALUSrc2_ID_0 & \input_b~2_combout )))) # (!\input_a~135_combout  & (ALUSrc2_ID_0 & ((\input_b~2_combout ))))

	.dataa(\input_a~135_combout ),
	.datab(\PR|ALUSrc2_ID [0]),
	.datac(\input_b~4_combout ),
	.datad(\input_b~2_combout ),
	.cin(gnd),
	.combout(\input_b~84_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~84 .lut_mask = 16'hECA0;
defparam \input_b~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \input_b~85 (
// Equation(s):
// \input_b~85_combout  = (\input_b~84_combout ) # ((Result_EX_0 & \input_b~1_combout ))

	.dataa(Result_EX_0),
	.datab(\input_b~1_combout ),
	.datac(gnd),
	.datad(\input_b~84_combout ),
	.cin(gnd),
	.combout(\input_b~85_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~85 .lut_mask = 16'hFF88;
defparam \input_b~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N28
cycloneive_lcell_comb \input_a~136 (
// Equation(s):
// \input_a~136_combout  = (src1_hazard_t & ((\input_a~141_combout ))) # (!src1_hazard_t & (ALUSrc1_ID_0))

	.dataa(\PR|ALUSrc1_ID [0]),
	.datab(gnd),
	.datac(\HZ|src1_hazard_t~1_combout ),
	.datad(\input_a~141_combout ),
	.cin(gnd),
	.combout(\input_a~136_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~136 .lut_mask = 16'hFA0A;
defparam \input_a~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N30
cycloneive_lcell_comb \input_a~137 (
// Equation(s):
// \input_a~137_combout  = (always03 & (Result_EX_0 & (\input_a~58_combout ))) # (!always03 & ((\input_a~136_combout ) # ((Result_EX_0 & \input_a~58_combout ))))

	.dataa(\HZ|always0~8_combout ),
	.datab(Result_EX_0),
	.datac(\input_a~58_combout ),
	.datad(\input_a~136_combout ),
	.cin(gnd),
	.combout(\input_a~137_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~137 .lut_mask = 16'hD5C0;
defparam \input_a~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N6
cycloneive_lcell_comb \halt_reg~10 (
// Equation(s):
// \halt_reg~10_combout  = (!ALUOP_ID_2 & !ALUOP_ID_3)

	.dataa(gnd),
	.datab(gnd),
	.datac(\PR|ALUOP_ID [2]),
	.datad(\PR|ALUOP_ID [3]),
	.cin(gnd),
	.combout(\halt_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~10 .lut_mask = 16'h000F;
defparam \halt_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \input_b~86 (
// Equation(s):
// \input_b~86_combout  = (\input_b~1_combout  & Result_EX_7)

	.dataa(gnd),
	.datab(gnd),
	.datac(\input_b~1_combout ),
	.datad(Result_EX_7),
	.cin(gnd),
	.combout(\input_b~86_combout ),
	.cout());
// synopsys translate_off
defparam \input_b~86 .lut_mask = 16'hF000;
defparam \input_b~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \input_a~138 (
// Equation(s):
// \input_a~138_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_3)) # (!MemToReg_MEM1 & ((CalcData_MEM_3)))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [3]),
	.datad(\PR|CalcData_MEM [3]),
	.cin(gnd),
	.combout(\input_a~138_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~138 .lut_mask = 16'hC480;
defparam \input_a~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \pc_next[3]~6 (
// Equation(s):
// \pc_next[3]~6_combout  = (\pc[22]~34_combout  & ((\input_a~138_combout ) # ((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & (((ALUSrc1_ID_3 & !\pc[22]~38_combout ))))

	.dataa(\input_a~138_combout ),
	.datab(\pc[22]~34_combout ),
	.datac(\PR|ALUSrc1_ID [3]),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~6 .lut_mask = 16'hCCB8;
defparam \pc_next[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \input_a~139 (
// Equation(s):
// \input_a~139_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_5)) # (!MemToReg_MEM1 & ((CalcData_MEM_5)))))

	.dataa(\PR|ReadData_MEM [5]),
	.datab(\PR|CalcData_MEM [5]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~139_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~139 .lut_mask = 16'hA0C0;
defparam \input_a~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \pc_next[5]~15 (
// Equation(s):
// \pc_next[5]~15_combout  = (\pc[22]~34_combout  & ((\input_a~139_combout ) # ((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & (((!\pc[22]~38_combout  & ALUSrc1_ID_5))))

	.dataa(\pc[22]~34_combout ),
	.datab(\input_a~139_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|ALUSrc1_ID [5]),
	.cin(gnd),
	.combout(\pc_next[5]~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~15 .lut_mask = 16'hADA8;
defparam \pc_next[5]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \pc_next[7]~23 (
// Equation(s):
// \pc_next[7]~23_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & ((\input_a~143_combout ))) # (!\pc[22]~34_combout  & (ALUSrc1_ID_7))))

	.dataa(\PR|ALUSrc1_ID [7]),
	.datab(\input_a~143_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[7]~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~23 .lut_mask = 16'hFC0A;
defparam \pc_next[7]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N14
cycloneive_lcell_comb \pc_next[6]~27 (
// Equation(s):
// \pc_next[6]~27_combout  = (\pc[22]~38_combout  & (((Instr_ID_4) # (\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_6 & ((!\pc[22]~34_combout ))))

	.dataa(\PR|ALUSrc1_ID [6]),
	.datab(\pc[22]~38_combout ),
	.datac(\PR|Instr_ID [4]),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~27 .lut_mask = 16'hCCE2;
defparam \pc_next[6]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N2
cycloneive_lcell_comb \pc_next[19]~71 (
// Equation(s):
// \pc_next[19]~71_combout  = (\pc[22]~34_combout  & ((\input_a~155_combout ) # ((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & (((ALUSrc1_ID_19 & !\pc[22]~38_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(\input_a~155_combout ),
	.datac(\PR|ALUSrc1_ID [19]),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[19]~71_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~71 .lut_mask = 16'hAAD8;
defparam \pc_next[19]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \pc_next[19]~72 (
// Equation(s):
// \pc_next[19]~72_combout  = (\pc_next[19]~71_combout  & (((Result_EX_19)) # (!\pc[22]~38_combout ))) # (!\pc_next[19]~71_combout  & (\pc[22]~38_combout  & ((Instr_ID_17))))

	.dataa(\pc_next[19]~71_combout ),
	.datab(\pc[22]~38_combout ),
	.datac(Result_EX_19),
	.datad(\PR|Instr_ID [17]),
	.cin(gnd),
	.combout(\pc_next[19]~72_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~72 .lut_mask = 16'hE6A2;
defparam \pc_next[19]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \pc_next[21]~79 (
// Equation(s):
// \pc_next[21]~79_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & (\input_a~157_combout )) # (!\pc[22]~34_combout  & ((ALUSrc1_ID_21)))))

	.dataa(\input_a~157_combout ),
	.datab(\PR|ALUSrc1_ID [21]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[21]~79_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~79 .lut_mask = 16'hFA0C;
defparam \pc_next[21]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \pc_next[21]~80 (
// Equation(s):
// \pc_next[21]~80_combout  = (\pc_next[21]~79_combout  & ((Result_EX_21) # ((!\pc[22]~38_combout )))) # (!\pc_next[21]~79_combout  & (((\pc[22]~38_combout  & Instr_ID_19))))

	.dataa(Result_EX_21),
	.datab(\pc_next[21]~79_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [19]),
	.cin(gnd),
	.combout(\pc_next[21]~80_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~80 .lut_mask = 16'hBC8C;
defparam \pc_next[21]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \pc_next[27]~103 (
// Equation(s):
// \pc_next[27]~103_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & (\input_a~163_combout )) # (!\pc[22]~34_combout  & ((ALUSrc1_ID_27)))))

	.dataa(\input_a~163_combout ),
	.datab(\PR|ALUSrc1_ID [27]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[27]~103_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~103 .lut_mask = 16'hFA0C;
defparam \pc_next[27]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N10
cycloneive_lcell_comb \pc[29]~29 (
// Equation(s):
// \pc[29]~29_combout  = (jump_ID_2 & (!jump_ID_1 & !jump_ID_0)) # (!jump_ID_2 & ((jump_ID_0)))

	.dataa(gnd),
	.datab(\PR|jump_ID [1]),
	.datac(\PR|jump_ID [2]),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\pc[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc[29]~29 .lut_mask = 16'h0F30;
defparam \pc[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N12
cycloneive_lcell_comb \pc_next[28]~114 (
// Equation(s):
// \pc_next[28]~114_combout  = (\pc[29]~30_combout  & (((\pc[29]~35_combout )))) # (!\pc[29]~30_combout  & ((\pc[29]~35_combout  & (ALUSrc1_ID_28)) # (!\pc[29]~35_combout  & ((\input_a~166_combout )))))

	.dataa(\pc[29]~30_combout ),
	.datab(\PR|ALUSrc1_ID [28]),
	.datac(\input_a~166_combout ),
	.datad(\pc[29]~35_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~114_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~114 .lut_mask = 16'hEE50;
defparam \pc_next[28]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N0
cycloneive_lcell_comb \Equal20~0 (
// Equation(s):
// \Equal20~0_combout  = (MemToReg_EX1 & (MemToReg_MEM1 & (src1_hazard_t & !always03)))

	.dataa(MemToReg_EX),
	.datab(\PR|MemToReg_MEM~q ),
	.datac(\HZ|src1_hazard_t~1_combout ),
	.datad(\HZ|always0~8_combout ),
	.cin(gnd),
	.combout(\Equal20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal20~0 .lut_mask = 16'h0080;
defparam \Equal20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!Selector141 & (!WideOr14 & ((Instr_IF_30) # (!WideOr211))))

	.dataa(\PR|Instr_IF [30]),
	.datab(\CU|WideOr21~2_combout ),
	.datac(\CU|Selector14~2_combout ),
	.datad(\CU|WideOr14~0_combout ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h000B;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (!Selector141 & ((Instr_IF_30) # (!WideOr211)))

	.dataa(gnd),
	.datab(\CU|Selector14~2_combout ),
	.datac(\CU|WideOr21~2_combout ),
	.datad(\PR|Instr_IF [30]),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h3303;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \input_ALUSrc2_ID~0 (
// Equation(s):
// \input_ALUSrc2_ID~0_combout  = (Selector141) # ((!Instr_IF_30 & (WideOr211 & !WideOr14)))

	.dataa(\PR|Instr_IF [30]),
	.datab(\CU|WideOr21~2_combout ),
	.datac(\CU|Selector14~2_combout ),
	.datad(\CU|WideOr14~0_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~0 .lut_mask = 16'hF0F4;
defparam \input_ALUSrc2_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \input_ALUSrc2_ID~1 (
// Equation(s):
// \input_ALUSrc2_ID~1_combout  = (Selector141) # ((WideOr14 & ((Instr_IF_30) # (!WideOr211))))

	.dataa(\PR|Instr_IF [30]),
	.datab(\CU|WideOr21~2_combout ),
	.datac(\CU|Selector14~2_combout ),
	.datad(\CU|WideOr14~0_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~1 .lut_mask = 16'hFBF0;
defparam \input_ALUSrc2_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \input_ALUSrc2_ID~2 (
// Equation(s):
// \input_ALUSrc2_ID~2_combout  = (\input_ALUSrc2_ID~1_combout  & (((Instr_IF_10) # (!\input_ALUSrc2_ID~0_combout )))) # (!\input_ALUSrc2_ID~1_combout  & (Instr_IF_4 & (\input_ALUSrc2_ID~0_combout )))

	.dataa(\input_ALUSrc2_ID~1_combout ),
	.datab(\PR|Instr_IF [4]),
	.datac(\input_ALUSrc2_ID~0_combout ),
	.datad(\PR|Instr_IF [10]),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~2 .lut_mask = 16'hEA4A;
defparam \input_ALUSrc2_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \input_ALUSrc2_ID~3 (
// Equation(s):
// \input_ALUSrc2_ID~3_combout  = (\Equal2~0_combout  & ((\input_ALUSrc2_ID~2_combout  & ((Instr_IF_4))) # (!\input_ALUSrc2_ID~2_combout  & (rfifrdat2_4)))) # (!\Equal2~0_combout  & (((\input_ALUSrc2_ID~2_combout ))))

	.dataa(\RF|rfif.rdat2[4]~587_combout ),
	.datab(\Equal2~0_combout ),
	.datac(\input_ALUSrc2_ID~2_combout ),
	.datad(\PR|Instr_IF [4]),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~3 .lut_mask = 16'hF838;
defparam \input_ALUSrc2_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \input_ALUSrc2_ID~4 (
// Equation(s):
// \input_ALUSrc2_ID~4_combout  = (\input_ALUSrc2_ID~1_combout  & ((Instr_IF_9) # ((!\input_ALUSrc2_ID~0_combout )))) # (!\input_ALUSrc2_ID~1_combout  & (((\input_ALUSrc2_ID~0_combout  & Instr_IF_3))))

	.dataa(\input_ALUSrc2_ID~1_combout ),
	.datab(\PR|Instr_IF [9]),
	.datac(\input_ALUSrc2_ID~0_combout ),
	.datad(\PR|Instr_IF [3]),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~4 .lut_mask = 16'hDA8A;
defparam \input_ALUSrc2_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \input_ALUSrc2_ID~5 (
// Equation(s):
// \input_ALUSrc2_ID~5_combout  = (\Equal2~0_combout  & ((\input_ALUSrc2_ID~4_combout  & (Instr_IF_3)) # (!\input_ALUSrc2_ID~4_combout  & ((rfifrdat2_3))))) # (!\Equal2~0_combout  & (((\input_ALUSrc2_ID~4_combout ))))

	.dataa(\PR|Instr_IF [3]),
	.datab(\Equal2~0_combout ),
	.datac(\input_ALUSrc2_ID~4_combout ),
	.datad(\RF|rfif.rdat2[3]~608_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~5 .lut_mask = 16'hBCB0;
defparam \input_ALUSrc2_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \input_ALUSrc2_ID~6 (
// Equation(s):
// \input_ALUSrc2_ID~6_combout  = (\input_ALUSrc2_ID~0_combout  & ((\input_ALUSrc2_ID~1_combout  & ((Instr_IF_8))) # (!\input_ALUSrc2_ID~1_combout  & (Instr_IF_2)))) # (!\input_ALUSrc2_ID~0_combout  & (((\input_ALUSrc2_ID~1_combout ))))

	.dataa(\input_ALUSrc2_ID~0_combout ),
	.datab(\PR|Instr_IF [2]),
	.datac(\PR|Instr_IF [8]),
	.datad(\input_ALUSrc2_ID~1_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~6 .lut_mask = 16'hF588;
defparam \input_ALUSrc2_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \input_ALUSrc2_ID~7 (
// Equation(s):
// \input_ALUSrc2_ID~7_combout  = (\input_ALUSrc2_ID~6_combout  & (((Instr_IF_2)) # (!\Equal2~0_combout ))) # (!\input_ALUSrc2_ID~6_combout  & (\Equal2~0_combout  & ((rfifrdat2_2))))

	.dataa(\input_ALUSrc2_ID~6_combout ),
	.datab(\Equal2~0_combout ),
	.datac(\PR|Instr_IF [2]),
	.datad(\RF|rfif.rdat2[2]~629_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~7 .lut_mask = 16'hE6A2;
defparam \input_ALUSrc2_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \input_ALUSrc2_ID~8 (
// Equation(s):
// \input_ALUSrc2_ID~8_combout  = (\input_ALUSrc2_ID~1_combout  & (((Instr_IF_7) # (!\input_ALUSrc2_ID~0_combout )))) # (!\input_ALUSrc2_ID~1_combout  & (Instr_IF_1 & (\input_ALUSrc2_ID~0_combout )))

	.dataa(\input_ALUSrc2_ID~1_combout ),
	.datab(\PR|Instr_IF [1]),
	.datac(\input_ALUSrc2_ID~0_combout ),
	.datad(\PR|Instr_IF [7]),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~8 .lut_mask = 16'hEA4A;
defparam \input_ALUSrc2_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \input_ALUSrc2_ID~9 (
// Equation(s):
// \input_ALUSrc2_ID~9_combout  = (\input_ALUSrc2_ID~8_combout  & ((Instr_IF_1) # ((!\Equal2~0_combout )))) # (!\input_ALUSrc2_ID~8_combout  & (((rfifrdat2_1 & \Equal2~0_combout ))))

	.dataa(\input_ALUSrc2_ID~8_combout ),
	.datab(\PR|Instr_IF [1]),
	.datac(\RF|rfif.rdat2[1]~650_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~9 .lut_mask = 16'hD8AA;
defparam \input_ALUSrc2_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \input_ALUSrc2_ID~10 (
// Equation(s):
// \input_ALUSrc2_ID~10_combout  = (\input_ALUSrc2_ID~0_combout  & ((\input_ALUSrc2_ID~1_combout  & (Instr_IF_6)) # (!\input_ALUSrc2_ID~1_combout  & ((Instr_IF_0))))) # (!\input_ALUSrc2_ID~0_combout  & (((\input_ALUSrc2_ID~1_combout ))))

	.dataa(\PR|Instr_IF [6]),
	.datab(\input_ALUSrc2_ID~0_combout ),
	.datac(\PR|Instr_IF [0]),
	.datad(\input_ALUSrc2_ID~1_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~10 .lut_mask = 16'hBBC0;
defparam \input_ALUSrc2_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \input_ALUSrc2_ID~11 (
// Equation(s):
// \input_ALUSrc2_ID~11_combout  = (\Equal2~0_combout  & ((\input_ALUSrc2_ID~10_combout  & (Instr_IF_0)) # (!\input_ALUSrc2_ID~10_combout  & ((rfifrdat2_0))))) # (!\Equal2~0_combout  & (((\input_ALUSrc2_ID~10_combout ))))

	.dataa(\PR|Instr_IF [0]),
	.datab(\Equal2~0_combout ),
	.datac(\RF|rfif.rdat2[0]~671_combout ),
	.datad(\input_ALUSrc2_ID~10_combout ),
	.cin(gnd),
	.combout(\input_ALUSrc2_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \input_ALUSrc2_ID~11 .lut_mask = 16'hBBC0;
defparam \input_ALUSrc2_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \Equal27~0 (
// Equation(s):
// \Equal27~0_combout  = (src2_hazard_t & (!always01 & ((!MemToReg_EX1) # (!MemToReg_MEM1))))

	.dataa(\HZ|src2_hazard_t~2_combout ),
	.datab(\HZ|always0~1_combout ),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(MemToReg_EX),
	.cin(gnd),
	.combout(\Equal27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal27~0 .lut_mask = 16'h0222;
defparam \Equal27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N18
cycloneive_lcell_comb \input_a~141 (
// Equation(s):
// \input_a~141_combout  = (MemToReg_MEM1 & (((ReadData_MEM_0 & !MemToReg_EX1)))) # (!MemToReg_MEM1 & (CalcData_MEM_0))

	.dataa(\PR|CalcData_MEM [0]),
	.datab(\PR|ReadData_MEM [0]),
	.datac(MemToReg_EX),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~141_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~141 .lut_mask = 16'h0CAA;
defparam \input_a~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \input_a~142 (
// Equation(s):
// \input_a~142_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_2))) # (!MemToReg_MEM1 & (CalcData_MEM_2))))

	.dataa(\PR|CalcData_MEM [2]),
	.datab(\PR|MemToReg_MEM~q ),
	.datac(\PR|ReadData_MEM [2]),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~142_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~142 .lut_mask = 16'hE200;
defparam \input_a~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \input_a~143 (
// Equation(s):
// \input_a~143_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_7)) # (!MemToReg_MEM1 & ((CalcData_MEM_7)))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|MemToReg_MEM~q ),
	.datac(\PR|ReadData_MEM [7]),
	.datad(\PR|CalcData_MEM [7]),
	.cin(gnd),
	.combout(\input_a~143_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~143 .lut_mask = 16'hA280;
defparam \input_a~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \input_a~145 (
// Equation(s):
// \input_a~145_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_9)) # (!MemToReg_MEM1 & ((CalcData_MEM_9)))))

	.dataa(\PR|ReadData_MEM [9]),
	.datab(\PR|CalcData_MEM [9]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~145_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~145 .lut_mask = 16'hA0C0;
defparam \input_a~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N6
cycloneive_lcell_comb \input_a~152 (
// Equation(s):
// \input_a~152_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_14))) # (!MemToReg_MEM1 & (CalcData_MEM_14))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|MemToReg_MEM~q ),
	.datac(\PR|CalcData_MEM [14]),
	.datad(\PR|ReadData_MEM [14]),
	.cin(gnd),
	.combout(\input_a~152_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~152 .lut_mask = 16'hA820;
defparam \input_a~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \input_a~155 (
// Equation(s):
// \input_a~155_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_19))) # (!MemToReg_MEM1 & (CalcData_MEM_19))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\Equal24~0_combout ),
	.datac(\PR|CalcData_MEM [19]),
	.datad(\PR|ReadData_MEM [19]),
	.cin(gnd),
	.combout(\input_a~155_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~155 .lut_mask = 16'hC840;
defparam \input_a~155 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \input_a~157 (
// Equation(s):
// \input_a~157_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_21)) # (!MemToReg_MEM1 & ((CalcData_MEM_21)))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [21]),
	.datad(\PR|CalcData_MEM [21]),
	.cin(gnd),
	.combout(\input_a~157_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~157 .lut_mask = 16'hC480;
defparam \input_a~157 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \input_a~162 (
// Equation(s):
// \input_a~162_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_24))) # (!MemToReg_MEM1 & (CalcData_MEM_24))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|CalcData_MEM [24]),
	.datac(\PR|ReadData_MEM [24]),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~162_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~162 .lut_mask = 16'hE400;
defparam \input_a~162 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \input_a~163 (
// Equation(s):
// \input_a~163_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_27))) # (!MemToReg_MEM1 & (CalcData_MEM_27))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|CalcData_MEM [27]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|ReadData_MEM [27]),
	.cin(gnd),
	.combout(\input_a~163_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~163 .lut_mask = 16'hE040;
defparam \input_a~163 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \input_a~165 (
// Equation(s):
// \input_a~165_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_29))) # (!MemToReg_MEM1 & (CalcData_MEM_29))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|CalcData_MEM [29]),
	.datac(\PR|ReadData_MEM [29]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~165_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~165 .lut_mask = 16'hA088;
defparam \input_a~165 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \input_a~166 (
// Equation(s):
// \input_a~166_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_28))) # (!MemToReg_MEM1 & (CalcData_MEM_28))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|CalcData_MEM [28]),
	.datac(\PR|ReadData_MEM [28]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~166_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~166 .lut_mask = 16'hA088;
defparam \input_a~166 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N9
dffeas \pc[1] (
	.clk(CLK),
	.d(\pc_next~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[1]~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_1),
	.prn(vcc));
// synopsys translate_off
defparam \pc[1] .is_wysiwyg = "true";
defparam \pc[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N29
dffeas \pc[0] (
	.clk(CLK),
	.d(\pc_next~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[1]~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_0),
	.prn(vcc));
// synopsys translate_off
defparam \pc[0] .is_wysiwyg = "true";
defparam \pc[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N5
dffeas \pc[3] (
	.clk(CLK),
	.d(\pc_next[3]~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_3),
	.prn(vcc));
// synopsys translate_off
defparam \pc[3] .is_wysiwyg = "true";
defparam \pc[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N9
dffeas \pc[2] (
	.clk(CLK),
	.d(\pc_next[2]~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_2),
	.prn(vcc));
// synopsys translate_off
defparam \pc[2] .is_wysiwyg = "true";
defparam \pc[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N17
dffeas \pc[5] (
	.clk(CLK),
	.d(\pc_next[5]~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_5),
	.prn(vcc));
// synopsys translate_off
defparam \pc[5] .is_wysiwyg = "true";
defparam \pc[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \pc[4] (
	.clk(CLK),
	.d(\pc_next[4]~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_4),
	.prn(vcc));
// synopsys translate_off
defparam \pc[4] .is_wysiwyg = "true";
defparam \pc[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N27
dffeas \pc[7] (
	.clk(CLK),
	.d(\pc_next[7]~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_7),
	.prn(vcc));
// synopsys translate_off
defparam \pc[7] .is_wysiwyg = "true";
defparam \pc[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N23
dffeas \pc[6] (
	.clk(CLK),
	.d(\pc_next[6]~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_6),
	.prn(vcc));
// synopsys translate_off
defparam \pc[6] .is_wysiwyg = "true";
defparam \pc[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N13
dffeas \pc[9] (
	.clk(CLK),
	.d(\pc_next[9]~34_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_9),
	.prn(vcc));
// synopsys translate_off
defparam \pc[9] .is_wysiwyg = "true";
defparam \pc[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \pc[8] (
	.clk(CLK),
	.d(\pc_next[8]~38_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_8),
	.prn(vcc));
// synopsys translate_off
defparam \pc[8] .is_wysiwyg = "true";
defparam \pc[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N25
dffeas \pc[11] (
	.clk(CLK),
	.d(\pc_next[11]~42_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_11),
	.prn(vcc));
// synopsys translate_off
defparam \pc[11] .is_wysiwyg = "true";
defparam \pc[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N29
dffeas \pc[10] (
	.clk(CLK),
	.d(\pc_next[10]~46_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_10),
	.prn(vcc));
// synopsys translate_off
defparam \pc[10] .is_wysiwyg = "true";
defparam \pc[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N9
dffeas \pc[13] (
	.clk(CLK),
	.d(\pc_next[13]~50_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_13),
	.prn(vcc));
// synopsys translate_off
defparam \pc[13] .is_wysiwyg = "true";
defparam \pc[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N5
dffeas \pc[12] (
	.clk(CLK),
	.d(\pc_next[12]~54_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_12),
	.prn(vcc));
// synopsys translate_off
defparam \pc[12] .is_wysiwyg = "true";
defparam \pc[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N27
dffeas \pc[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_next[15]~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_15),
	.prn(vcc));
// synopsys translate_off
defparam \pc[15] .is_wysiwyg = "true";
defparam \pc[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N1
dffeas \pc[14] (
	.clk(CLK),
	.d(\pc_next[14]~62_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_14),
	.prn(vcc));
// synopsys translate_off
defparam \pc[14] .is_wysiwyg = "true";
defparam \pc[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N21
dffeas \pc[17] (
	.clk(CLK),
	.d(\pc_next[17]~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_17),
	.prn(vcc));
// synopsys translate_off
defparam \pc[17] .is_wysiwyg = "true";
defparam \pc[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N13
dffeas \pc[16] (
	.clk(CLK),
	.d(\pc_next[16]~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_16),
	.prn(vcc));
// synopsys translate_off
defparam \pc[16] .is_wysiwyg = "true";
defparam \pc[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N25
dffeas \pc[19] (
	.clk(CLK),
	.d(\pc_next[19]~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_19),
	.prn(vcc));
// synopsys translate_off
defparam \pc[19] .is_wysiwyg = "true";
defparam \pc[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N5
dffeas \pc[18] (
	.clk(CLK),
	.d(\pc_next[18]~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_18),
	.prn(vcc));
// synopsys translate_off
defparam \pc[18] .is_wysiwyg = "true";
defparam \pc[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N21
dffeas \pc[21] (
	.clk(CLK),
	.d(\pc_next[21]~82_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_21),
	.prn(vcc));
// synopsys translate_off
defparam \pc[21] .is_wysiwyg = "true";
defparam \pc[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N19
dffeas \pc[20] (
	.clk(CLK),
	.d(\pc_next[20]~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_20),
	.prn(vcc));
// synopsys translate_off
defparam \pc[20] .is_wysiwyg = "true";
defparam \pc[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N13
dffeas \pc[23] (
	.clk(CLK),
	.d(\pc_next[23]~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_23),
	.prn(vcc));
// synopsys translate_off
defparam \pc[23] .is_wysiwyg = "true";
defparam \pc[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N15
dffeas \pc[22] (
	.clk(CLK),
	.d(\pc_next[22]~94_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_22),
	.prn(vcc));
// synopsys translate_off
defparam \pc[22] .is_wysiwyg = "true";
defparam \pc[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N9
dffeas \pc[25] (
	.clk(CLK),
	.d(\pc_next[25]~98_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_25),
	.prn(vcc));
// synopsys translate_off
defparam \pc[25] .is_wysiwyg = "true";
defparam \pc[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \pc[24] (
	.clk(CLK),
	.d(\pc_next[24]~102_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_24),
	.prn(vcc));
// synopsys translate_off
defparam \pc[24] .is_wysiwyg = "true";
defparam \pc[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N15
dffeas \pc[27] (
	.clk(CLK),
	.d(\pc_next[27]~106_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_27),
	.prn(vcc));
// synopsys translate_off
defparam \pc[27] .is_wysiwyg = "true";
defparam \pc[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N19
dffeas \pc[26] (
	.clk(CLK),
	.d(\pc_next[26]~110_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC_enable~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_26),
	.prn(vcc));
// synopsys translate_off
defparam \pc[26] .is_wysiwyg = "true";
defparam \pc[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N25
dffeas \pc[29] (
	.clk(CLK),
	.d(\pc_next[29]~113_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_29),
	.prn(vcc));
// synopsys translate_off
defparam \pc[29] .is_wysiwyg = "true";
defparam \pc[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N3
dffeas \pc[28] (
	.clk(CLK),
	.d(\pc_next[28]~116_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_28),
	.prn(vcc));
// synopsys translate_off
defparam \pc[28] .is_wysiwyg = "true";
defparam \pc[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N5
dffeas \pc[31] (
	.clk(CLK),
	.d(\pc_next[31]~119_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_31),
	.prn(vcc));
// synopsys translate_off
defparam \pc[31] .is_wysiwyg = "true";
defparam \pc[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N11
dffeas \pc[30] (
	.clk(CLK),
	.d(\pc_next[30]~122_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[31]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_30),
	.prn(vcc));
// synopsys translate_off
defparam \pc[30] .is_wysiwyg = "true";
defparam \pc[30] .power_up = "low";
// synopsys translate_on

// Location: DDIOOUTCELL_X47_Y0_N11
dffeas halt_reg(
	.clk(!CLK),
	.d(\halt_reg~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(halt_reg1),
	.prn(vcc));
// synopsys translate_off
defparam halt_reg.is_wysiwyg = "true";
defparam halt_reg.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \Equal8~0 (
// Equation(s):
// \Equal8~0_combout  = (!jump_ID_1 & (!jump_ID_2 & jump_ID_0))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(gnd),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal8~0 .lut_mask = 16'h1100;
defparam \Equal8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Equal24~0 (
// Equation(s):
// \Equal24~0_combout  = (!always03 & (src1_hazard_t & ((!MemToReg_EX1) # (!MemToReg_MEM1))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(MemToReg_EX),
	.datac(\HZ|always0~8_combout ),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\Equal24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal24~0 .lut_mask = 16'h0700;
defparam \Equal24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \Equal8~1 (
// Equation(s):
// \Equal8~1_combout  = (jump_ID_1 & (!jump_ID_2 & !jump_ID_0))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(gnd),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\Equal8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal8~1 .lut_mask = 16'h0022;
defparam \Equal8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \pc[0]~37 (
// Equation(s):
// \pc[0]~37_combout  = (\Equal8~1_combout  & ((always03 & (!MemToReg_EX1)) # (!always03 & ((!src1_hazard_t)))))

	.dataa(MemToReg_EX),
	.datab(\Equal8~1_combout ),
	.datac(\HZ|always0~8_combout ),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\pc[0]~37_combout ),
	.cout());
// synopsys translate_off
defparam \pc[0]~37 .lut_mask = 16'h404C;
defparam \pc[0]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \pc_next~0 (
// Equation(s):
// \pc_next~0_combout  = (\pc[0]~33_combout  & ((\pc[0]~37_combout  & ((ALUSrc1_ID_1))) # (!\pc[0]~37_combout  & (nextPC_ID_1)))) # (!\pc[0]~33_combout  & (\pc[0]~37_combout ))

	.dataa(\pc[0]~33_combout ),
	.datab(\pc[0]~37_combout ),
	.datac(\PR|nextPC_ID [1]),
	.datad(\PR|ALUSrc1_ID [1]),
	.cin(gnd),
	.combout(\pc_next~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~0 .lut_mask = 16'hEC64;
defparam \pc_next~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \input_a~132 (
// Equation(s):
// \input_a~132_combout  = (MemToReg_MEM1 & (ReadData_MEM_1)) # (!MemToReg_MEM1 & ((CalcData_MEM_1)))

	.dataa(gnd),
	.datab(\PR|ReadData_MEM [1]),
	.datac(\PR|CalcData_MEM [1]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~132_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~132 .lut_mask = 16'hCCF0;
defparam \input_a~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \Equal22~0 (
// Equation(s):
// \Equal22~0_combout  = (always03) # (src1_hazard_t)

	.dataa(gnd),
	.datab(gnd),
	.datac(\HZ|always0~8_combout ),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\Equal22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal22~0 .lut_mask = 16'hFFF0;
defparam \Equal22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \pc[0]~25 (
// Equation(s):
// \pc[0]~25_combout  = (jump_ID_1 & (!jump_ID_2 & (\Equal22~0_combout  & !jump_ID_0)))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(\Equal22~0_combout ),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\pc[0]~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc[0]~25 .lut_mask = 16'h0020;
defparam \pc[0]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \pc_next~1 (
// Equation(s):
// \pc_next~1_combout  = (\pc[0]~25_combout  & ((\pc_next~0_combout  & (!Result_EX_1)) # (!\pc_next~0_combout  & ((\input_a~132_combout )))))

	.dataa(\pc_next~0_combout ),
	.datab(Result_EX_1),
	.datac(\input_a~132_combout ),
	.datad(\pc[0]~25_combout ),
	.cin(gnd),
	.combout(\pc_next~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~1 .lut_mask = 16'h7200;
defparam \pc_next~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \pc_next~2 (
// Equation(s):
// \pc_next~2_combout  = (!\Equal8~0_combout  & ((\pc_next~0_combout  & ((!\pc_next~1_combout ))) # (!\pc_next~0_combout  & (\Equal24~0_combout  & \pc_next~1_combout ))))

	.dataa(\Equal8~0_combout ),
	.datab(\Equal24~0_combout ),
	.datac(\pc_next~0_combout ),
	.datad(\pc_next~1_combout ),
	.cin(gnd),
	.combout(\pc_next~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~2 .lut_mask = 16'h0450;
defparam \pc_next~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N26
cycloneive_lcell_comb \branch~0 (
// Equation(s):
// \branch~0_combout  = (jump_ID_1 & (!jump_ID_2 & ((Equal11) # (!jump_ID_0)))) # (!jump_ID_1 & ((jump_ID_2 & (!jump_ID_0 & !Equal11)) # (!jump_ID_2 & (jump_ID_0))))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(\PR|jump_ID [0]),
	.datad(\ALU|Equal11~11_combout ),
	.cin(gnd),
	.combout(\branch~0_combout ),
	.cout());
// synopsys translate_off
defparam \branch~0 .lut_mask = 16'h3216;
defparam \branch~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \pc[1]~26 (
// Equation(s):
// \pc[1]~26_combout  = (Equal11 & ((jump_ID_1) # ((jump_ID_0)))) # (!Equal11 & ((jump_ID_2) # (jump_ID_1 $ (jump_ID_0))))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(\PR|jump_ID [0]),
	.datad(\ALU|Equal11~11_combout ),
	.cin(gnd),
	.combout(\pc[1]~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc[1]~26 .lut_mask = 16'hFADE;
defparam \pc[1]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \pc[1]~27 (
// Equation(s):
// \pc[1]~27_combout  = (always1 & (\pc[1]~26_combout  & ((\branch~0_combout ) # (!always0))))

	.dataa(always1),
	.datab(always0),
	.datac(\branch~0_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc[1]~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc[1]~27 .lut_mask = 16'hA200;
defparam \pc[1]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \pc[0]~24 (
// Equation(s):
// \pc[0]~24_combout  = jump_ID_2 $ (((jump_ID_1) # (jump_ID_0)))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(gnd),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\pc[0]~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc[0]~24 .lut_mask = 16'h3366;
defparam \pc[0]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N0
cycloneive_lcell_comb \pc[0]~33 (
// Equation(s):
// \pc[0]~33_combout  = (\Equal8~1_combout  & (!always03 & ((!src1_hazard_t)))) # (!\Equal8~1_combout  & (((\pc[0]~24_combout ))))

	.dataa(\HZ|always0~8_combout ),
	.datab(\pc[0]~24_combout ),
	.datac(\Equal8~1_combout ),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\pc[0]~33_combout ),
	.cout());
// synopsys translate_off
defparam \pc[0]~33 .lut_mask = 16'h0C5C;
defparam \pc[0]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \pc_next~3 (
// Equation(s):
// \pc_next~3_combout  = (\pc[0]~33_combout  & ((\pc[0]~37_combout  & ((ALUSrc1_ID_0))) # (!\pc[0]~37_combout  & (nextPC_ID_0)))) # (!\pc[0]~33_combout  & (((\pc[0]~37_combout ))))

	.dataa(\PR|nextPC_ID [0]),
	.datab(\pc[0]~33_combout ),
	.datac(\pc[0]~37_combout ),
	.datad(\PR|ALUSrc1_ID [0]),
	.cin(gnd),
	.combout(\pc_next~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~3 .lut_mask = 16'hF838;
defparam \pc_next~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N8
cycloneive_lcell_comb \input_a~135 (
// Equation(s):
// \input_a~135_combout  = (MemToReg_MEM1 & ((ReadData_MEM_0))) # (!MemToReg_MEM1 & (CalcData_MEM_0))

	.dataa(\PR|CalcData_MEM [0]),
	.datab(\PR|ReadData_MEM [0]),
	.datac(gnd),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~135_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~135 .lut_mask = 16'hCCAA;
defparam \input_a~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \pc_next~4 (
// Equation(s):
// \pc_next~4_combout  = (\pc[0]~25_combout  & ((\pc_next~3_combout  & (!Result_EX_0)) # (!\pc_next~3_combout  & ((\input_a~135_combout )))))

	.dataa(Result_EX_0),
	.datab(\pc_next~3_combout ),
	.datac(\input_a~135_combout ),
	.datad(\pc[0]~25_combout ),
	.cin(gnd),
	.combout(\pc_next~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~4 .lut_mask = 16'h7400;
defparam \pc_next~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \pc_next~5 (
// Equation(s):
// \pc_next~5_combout  = (!\Equal8~0_combout  & ((\pc_next~4_combout  & (\Equal24~0_combout  & !\pc_next~3_combout )) # (!\pc_next~4_combout  & ((\pc_next~3_combout )))))

	.dataa(\Equal8~0_combout ),
	.datab(\pc_next~4_combout ),
	.datac(\Equal24~0_combout ),
	.datad(\pc_next~3_combout ),
	.cin(gnd),
	.combout(\pc_next~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~5 .lut_mask = 16'h1140;
defparam \pc_next~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \pc_next_plus4[2]~0 (
// Equation(s):
// \pc_next_plus4[2]~0_combout  = pc_2 $ (VCC)
// \pc_next_plus4[2]~1  = CARRY(pc_2)

	.dataa(gnd),
	.datab(pc_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pc_next_plus4[2]~0_combout ),
	.cout(\pc_next_plus4[2]~1 ));
// synopsys translate_off
defparam \pc_next_plus4[2]~0 .lut_mask = 16'h33CC;
defparam \pc_next_plus4[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \pc_next_plus4[3]~2 (
// Equation(s):
// \pc_next_plus4[3]~2_combout  = (pc_3 & (!\pc_next_plus4[2]~1 )) # (!pc_3 & ((\pc_next_plus4[2]~1 ) # (GND)))
// \pc_next_plus4[3]~3  = CARRY((!\pc_next_plus4[2]~1 ) # (!pc_3))

	.dataa(gnd),
	.datab(pc_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[2]~1 ),
	.combout(\pc_next_plus4[3]~2_combout ),
	.cout(\pc_next_plus4[3]~3 ));
// synopsys translate_off
defparam \pc_next_plus4[3]~2 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \pc_next_branch[3]~2 (
// Equation(s):
// \pc_next_branch[3]~2_combout  = (Instr_ID_1 & ((nextPC_ID_3 & (\pc_next_branch[2]~1  & VCC)) # (!nextPC_ID_3 & (!\pc_next_branch[2]~1 )))) # (!Instr_ID_1 & ((nextPC_ID_3 & (!\pc_next_branch[2]~1 )) # (!nextPC_ID_3 & ((\pc_next_branch[2]~1 ) # (GND)))))
// \pc_next_branch[3]~3  = CARRY((Instr_ID_1 & (!nextPC_ID_3 & !\pc_next_branch[2]~1 )) # (!Instr_ID_1 & ((!\pc_next_branch[2]~1 ) # (!nextPC_ID_3))))

	.dataa(\PR|Instr_ID [1]),
	.datab(\PR|nextPC_ID [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[2]~1 ),
	.combout(\pc_next_branch[3]~2_combout ),
	.cout(\pc_next_branch[3]~3 ));
// synopsys translate_off
defparam \pc_next_branch[3]~2 .lut_mask = 16'h9617;
defparam \pc_next_branch[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N22
cycloneive_lcell_comb \pc[22]~38 (
// Equation(s):
// \pc[22]~38_combout  = (jump_ID_0) # ((always03 & !MemToReg_EX1))

	.dataa(\HZ|always0~8_combout ),
	.datab(MemToReg_EX),
	.datac(gnd),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\pc[22]~38_combout ),
	.cout());
// synopsys translate_off
defparam \pc[22]~38 .lut_mask = 16'hFF22;
defparam \pc[22]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \pc_next[3]~7 (
// Equation(s):
// \pc_next[3]~7_combout  = (\pc_next[3]~6_combout  & (((Result_EX_3) # (!\pc[22]~38_combout )))) # (!\pc_next[3]~6_combout  & (Instr_ID_1 & (\pc[22]~38_combout )))

	.dataa(\pc_next[3]~6_combout ),
	.datab(\PR|Instr_ID [1]),
	.datac(\pc[22]~38_combout ),
	.datad(Result_EX_3),
	.cin(gnd),
	.combout(\pc_next[3]~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~7 .lut_mask = 16'hEA4A;
defparam \pc_next[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N0
cycloneive_lcell_comb \pc[22]~28 (
// Equation(s):
// \pc[22]~28_combout  = (jump_ID_1 & (!jump_ID_2 & jump_ID_0)) # (!jump_ID_1 & (jump_ID_2 & !jump_ID_0))

	.dataa(gnd),
	.datab(\PR|jump_ID [1]),
	.datac(\PR|jump_ID [2]),
	.datad(\PR|jump_ID [0]),
	.cin(gnd),
	.combout(\pc[22]~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc[22]~28 .lut_mask = 16'h0C30;
defparam \pc[22]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \pc_next[3]~8 (
// Equation(s):
// \pc_next[3]~8_combout  = (\pc[22]~28_combout  & (\pc_next_branch[3]~2_combout )) # (!\pc[22]~28_combout  & ((\pc_next[3]~7_combout )))

	.dataa(gnd),
	.datab(\pc_next_branch[3]~2_combout ),
	.datac(\pc_next[3]~7_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~8 .lut_mask = 16'hCCF0;
defparam \pc_next[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \pc_next[27]~9 (
// Equation(s):
// \pc_next[27]~9_combout  = (jump_ID_1 & ((jump_ID_2) # ((jump_ID_0 & !Equal11)))) # (!jump_ID_1 & ((jump_ID_2 & ((jump_ID_0) # (Equal11))) # (!jump_ID_2 & (!jump_ID_0))))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(\PR|jump_ID [0]),
	.datad(\ALU|Equal11~11_combout ),
	.cin(gnd),
	.combout(\pc_next[27]~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~9 .lut_mask = 16'hCDE9;
defparam \pc_next[27]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \pc_next[3]~10 (
// Equation(s):
// \pc_next[3]~10_combout  = (\pc_next_plus4[3]~2_combout  & (((\pc_next[3]~8_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[3]~2_combout  & (\pc_next[3]~8_combout  & ((!\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[3]~2_combout ),
	.datab(\pc_next[3]~8_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[3]~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~10 .lut_mask = 16'h0ACE;
defparam \pc_next[3]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N20
cycloneive_lcell_comb \PC_enable~2 (
// Equation(s):
// \PC_enable~2_combout  = (always1 & ((\branch~0_combout ) # ((!MemToReg_EX1 & !Memwrite_EX1))))

	.dataa(always1),
	.datab(MemToReg_EX),
	.datac(Memwrite_EX),
	.datad(\branch~0_combout ),
	.cin(gnd),
	.combout(\PC_enable~2_combout ),
	.cout());
// synopsys translate_off
defparam \PC_enable~2 .lut_mask = 16'hAA02;
defparam \PC_enable~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \pc[22]~34 (
// Equation(s):
// \pc[22]~34_combout  = (!jump_ID_0 & ((always03) # (src1_hazard_t)))

	.dataa(\HZ|always0~8_combout ),
	.datab(\PR|jump_ID [0]),
	.datac(gnd),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\pc[22]~34_combout ),
	.cout());
// synopsys translate_off
defparam \pc[22]~34 .lut_mask = 16'h3322;
defparam \pc[22]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \pc_next[2]~11 (
// Equation(s):
// \pc_next[2]~11_combout  = (\pc[22]~38_combout  & (((Instr_ID_0) # (\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_2 & ((!\pc[22]~34_combout ))))

	.dataa(\pc[22]~38_combout ),
	.datab(\PR|ALUSrc1_ID [2]),
	.datac(\PR|Instr_ID [0]),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[2]~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~11 .lut_mask = 16'hAAE4;
defparam \pc_next[2]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \pc_next[2]~12 (
// Equation(s):
// \pc_next[2]~12_combout  = (\pc[22]~34_combout  & ((\pc_next[2]~11_combout  & ((Result_EX_2))) # (!\pc_next[2]~11_combout  & (\input_a~142_combout )))) # (!\pc[22]~34_combout  & (((\pc_next[2]~11_combout ))))

	.dataa(\input_a~142_combout ),
	.datab(\pc[22]~34_combout ),
	.datac(\pc_next[2]~11_combout ),
	.datad(Result_EX_2),
	.cin(gnd),
	.combout(\pc_next[2]~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~12 .lut_mask = 16'hF838;
defparam \pc_next[2]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \pc_next[2]~13 (
// Equation(s):
// \pc_next[2]~13_combout  = (\pc[22]~28_combout  & (\pc_next_branch[2]~0_combout )) # (!\pc[22]~28_combout  & ((\pc_next[2]~12_combout )))

	.dataa(\pc_next_branch[2]~0_combout ),
	.datab(\pc_next[2]~12_combout ),
	.datac(gnd),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[2]~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~13 .lut_mask = 16'hAACC;
defparam \pc_next[2]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \pc_next[2]~14 (
// Equation(s):
// \pc_next[2]~14_combout  = (\pc_next[2]~13_combout  & (((\pc_next_plus4[2]~0_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[2]~13_combout  & (\pc_next_plus4[2]~0_combout  & (!\pc[1]~26_combout )))

	.dataa(\pc_next[2]~13_combout ),
	.datab(\pc_next_plus4[2]~0_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[2]~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~14 .lut_mask = 16'h0CAE;
defparam \pc_next[2]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \pc_next_plus4[4]~4 (
// Equation(s):
// \pc_next_plus4[4]~4_combout  = (pc_4 & (\pc_next_plus4[3]~3  $ (GND))) # (!pc_4 & (!\pc_next_plus4[3]~3  & VCC))
// \pc_next_plus4[4]~5  = CARRY((pc_4 & !\pc_next_plus4[3]~3 ))

	.dataa(pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[3]~3 ),
	.combout(\pc_next_plus4[4]~4_combout ),
	.cout(\pc_next_plus4[4]~5 ));
// synopsys translate_off
defparam \pc_next_plus4[4]~4 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \pc_next_plus4[5]~6 (
// Equation(s):
// \pc_next_plus4[5]~6_combout  = (pc_5 & (!\pc_next_plus4[4]~5 )) # (!pc_5 & ((\pc_next_plus4[4]~5 ) # (GND)))
// \pc_next_plus4[5]~7  = CARRY((!\pc_next_plus4[4]~5 ) # (!pc_5))

	.dataa(gnd),
	.datab(pc_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[4]~5 ),
	.combout(\pc_next_plus4[5]~6_combout ),
	.cout(\pc_next_plus4[5]~7 ));
// synopsys translate_off
defparam \pc_next_plus4[5]~6 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \pc_next[5]~16 (
// Equation(s):
// \pc_next[5]~16_combout  = (\pc_next[5]~15_combout  & ((Result_EX_5) # ((!\pc[22]~38_combout )))) # (!\pc_next[5]~15_combout  & (((\pc[22]~38_combout  & Instr_ID_3))))

	.dataa(\pc_next[5]~15_combout ),
	.datab(Result_EX_5),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [3]),
	.cin(gnd),
	.combout(\pc_next[5]~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~16 .lut_mask = 16'hDA8A;
defparam \pc_next[5]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \pc_next_branch[4]~4 (
// Equation(s):
// \pc_next_branch[4]~4_combout  = ((Instr_ID_2 $ (nextPC_ID_4 $ (!\pc_next_branch[3]~3 )))) # (GND)
// \pc_next_branch[4]~5  = CARRY((Instr_ID_2 & ((nextPC_ID_4) # (!\pc_next_branch[3]~3 ))) # (!Instr_ID_2 & (nextPC_ID_4 & !\pc_next_branch[3]~3 )))

	.dataa(\PR|Instr_ID [2]),
	.datab(\PR|nextPC_ID [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[3]~3 ),
	.combout(\pc_next_branch[4]~4_combout ),
	.cout(\pc_next_branch[4]~5 ));
// synopsys translate_off
defparam \pc_next_branch[4]~4 .lut_mask = 16'h698E;
defparam \pc_next_branch[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \pc_next_branch[5]~6 (
// Equation(s):
// \pc_next_branch[5]~6_combout  = (nextPC_ID_5 & ((Instr_ID_3 & (\pc_next_branch[4]~5  & VCC)) # (!Instr_ID_3 & (!\pc_next_branch[4]~5 )))) # (!nextPC_ID_5 & ((Instr_ID_3 & (!\pc_next_branch[4]~5 )) # (!Instr_ID_3 & ((\pc_next_branch[4]~5 ) # (GND)))))
// \pc_next_branch[5]~7  = CARRY((nextPC_ID_5 & (!Instr_ID_3 & !\pc_next_branch[4]~5 )) # (!nextPC_ID_5 & ((!\pc_next_branch[4]~5 ) # (!Instr_ID_3))))

	.dataa(\PR|nextPC_ID [5]),
	.datab(\PR|Instr_ID [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[4]~5 ),
	.combout(\pc_next_branch[5]~6_combout ),
	.cout(\pc_next_branch[5]~7 ));
// synopsys translate_off
defparam \pc_next_branch[5]~6 .lut_mask = 16'h9617;
defparam \pc_next_branch[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \pc_next[5]~17 (
// Equation(s):
// \pc_next[5]~17_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[5]~6_combout ))) # (!\pc[22]~28_combout  & (\pc_next[5]~16_combout ))

	.dataa(\pc[22]~28_combout ),
	.datab(\pc_next[5]~16_combout ),
	.datac(\pc_next_branch[5]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_next[5]~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~17 .lut_mask = 16'hE4E4;
defparam \pc_next[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \pc_next[5]~18 (
// Equation(s):
// \pc_next[5]~18_combout  = (\pc_next_plus4[5]~6_combout  & (((\pc_next[5]~17_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[5]~6_combout  & (\pc_next[5]~17_combout  & ((!\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[5]~6_combout ),
	.datab(\pc_next[5]~17_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[5]~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~18 .lut_mask = 16'h0ACE;
defparam \pc_next[5]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N22
cycloneive_lcell_comb \input_a~140 (
// Equation(s):
// \input_a~140_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_4))) # (!MemToReg_MEM1 & (CalcData_MEM_4))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\Equal24~0_combout ),
	.datac(\PR|CalcData_MEM [4]),
	.datad(\PR|ReadData_MEM [4]),
	.cin(gnd),
	.combout(\input_a~140_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~140 .lut_mask = 16'hC840;
defparam \input_a~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N26
cycloneive_lcell_comb \pc_next[4]~19 (
// Equation(s):
// \pc_next[4]~19_combout  = (\pc[22]~38_combout  & ((Instr_ID_2) # ((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (((ALUSrc1_ID_4 & !\pc[22]~34_combout ))))

	.dataa(\PR|Instr_ID [2]),
	.datab(\pc[22]~38_combout ),
	.datac(\PR|ALUSrc1_ID [4]),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[4]~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~19 .lut_mask = 16'hCCB8;
defparam \pc_next[4]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N4
cycloneive_lcell_comb \pc_next[4]~20 (
// Equation(s):
// \pc_next[4]~20_combout  = (\pc[22]~34_combout  & ((\pc_next[4]~19_combout  & ((Result_EX_4))) # (!\pc_next[4]~19_combout  & (\input_a~140_combout )))) # (!\pc[22]~34_combout  & (((\pc_next[4]~19_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(\input_a~140_combout ),
	.datac(\pc_next[4]~19_combout ),
	.datad(Result_EX_4),
	.cin(gnd),
	.combout(\pc_next[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~20 .lut_mask = 16'hF858;
defparam \pc_next[4]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N22
cycloneive_lcell_comb \pc_next[4]~21 (
// Equation(s):
// \pc_next[4]~21_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[4]~4_combout ))) # (!\pc[22]~28_combout  & (\pc_next[4]~20_combout ))

	.dataa(gnd),
	.datab(\pc_next[4]~20_combout ),
	.datac(\pc_next_branch[4]~4_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[4]~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~21 .lut_mask = 16'hF0CC;
defparam \pc_next[4]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \pc_next[4]~22 (
// Equation(s):
// \pc_next[4]~22_combout  = (\pc_next_plus4[4]~4_combout  & (((\pc_next[4]~21_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[4]~4_combout  & (\pc_next[4]~21_combout  & ((!\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[4]~4_combout ),
	.datab(\pc_next[4]~21_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[4]~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~22 .lut_mask = 16'h0ACE;
defparam \pc_next[4]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \pc_next_branch[6]~8 (
// Equation(s):
// \pc_next_branch[6]~8_combout  = ((nextPC_ID_6 $ (Instr_ID_4 $ (!\pc_next_branch[5]~7 )))) # (GND)
// \pc_next_branch[6]~9  = CARRY((nextPC_ID_6 & ((Instr_ID_4) # (!\pc_next_branch[5]~7 ))) # (!nextPC_ID_6 & (Instr_ID_4 & !\pc_next_branch[5]~7 )))

	.dataa(\PR|nextPC_ID [6]),
	.datab(\PR|Instr_ID [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[5]~7 ),
	.combout(\pc_next_branch[6]~8_combout ),
	.cout(\pc_next_branch[6]~9 ));
// synopsys translate_off
defparam \pc_next_branch[6]~8 .lut_mask = 16'h698E;
defparam \pc_next_branch[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \pc_next_branch[7]~10 (
// Equation(s):
// \pc_next_branch[7]~10_combout  = (nextPC_ID_7 & ((Instr_ID_5 & (\pc_next_branch[6]~9  & VCC)) # (!Instr_ID_5 & (!\pc_next_branch[6]~9 )))) # (!nextPC_ID_7 & ((Instr_ID_5 & (!\pc_next_branch[6]~9 )) # (!Instr_ID_5 & ((\pc_next_branch[6]~9 ) # (GND)))))
// \pc_next_branch[7]~11  = CARRY((nextPC_ID_7 & (!Instr_ID_5 & !\pc_next_branch[6]~9 )) # (!nextPC_ID_7 & ((!\pc_next_branch[6]~9 ) # (!Instr_ID_5))))

	.dataa(\PR|nextPC_ID [7]),
	.datab(\PR|Instr_ID [5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[6]~9 ),
	.combout(\pc_next_branch[7]~10_combout ),
	.cout(\pc_next_branch[7]~11 ));
// synopsys translate_off
defparam \pc_next_branch[7]~10 .lut_mask = 16'h9617;
defparam \pc_next_branch[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \pc_next[7]~24 (
// Equation(s):
// \pc_next[7]~24_combout  = (\pc_next[7]~23_combout  & ((Result_EX_7) # ((!\pc[22]~38_combout )))) # (!\pc_next[7]~23_combout  & (((\pc[22]~38_combout  & Instr_ID_5))))

	.dataa(\pc_next[7]~23_combout ),
	.datab(Result_EX_7),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [5]),
	.cin(gnd),
	.combout(\pc_next[7]~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~24 .lut_mask = 16'hDA8A;
defparam \pc_next[7]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N28
cycloneive_lcell_comb \pc_next[7]~25 (
// Equation(s):
// \pc_next[7]~25_combout  = (\pc[22]~28_combout  & (\pc_next_branch[7]~10_combout )) # (!\pc[22]~28_combout  & ((\pc_next[7]~24_combout )))

	.dataa(\pc[22]~28_combout ),
	.datab(gnd),
	.datac(\pc_next_branch[7]~10_combout ),
	.datad(\pc_next[7]~24_combout ),
	.cin(gnd),
	.combout(\pc_next[7]~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~25 .lut_mask = 16'hF5A0;
defparam \pc_next[7]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \pc_next_plus4[6]~8 (
// Equation(s):
// \pc_next_plus4[6]~8_combout  = (pc_6 & (\pc_next_plus4[5]~7  $ (GND))) # (!pc_6 & (!\pc_next_plus4[5]~7  & VCC))
// \pc_next_plus4[6]~9  = CARRY((pc_6 & !\pc_next_plus4[5]~7 ))

	.dataa(pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[5]~7 ),
	.combout(\pc_next_plus4[6]~8_combout ),
	.cout(\pc_next_plus4[6]~9 ));
// synopsys translate_off
defparam \pc_next_plus4[6]~8 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \pc_next_plus4[7]~10 (
// Equation(s):
// \pc_next_plus4[7]~10_combout  = (pc_7 & (!\pc_next_plus4[6]~9 )) # (!pc_7 & ((\pc_next_plus4[6]~9 ) # (GND)))
// \pc_next_plus4[7]~11  = CARRY((!\pc_next_plus4[6]~9 ) # (!pc_7))

	.dataa(gnd),
	.datab(pc_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[6]~9 ),
	.combout(\pc_next_plus4[7]~10_combout ),
	.cout(\pc_next_plus4[7]~11 ));
// synopsys translate_off
defparam \pc_next_plus4[7]~10 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \pc_next[7]~26 (
// Equation(s):
// \pc_next[7]~26_combout  = (\pc_next[7]~25_combout  & (((\pc_next_plus4[7]~10_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[7]~25_combout  & (\pc_next_plus4[7]~10_combout  & (!\pc[1]~26_combout )))

	.dataa(\pc_next[7]~25_combout ),
	.datab(\pc_next_plus4[7]~10_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[7]~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~26 .lut_mask = 16'h0CAE;
defparam \pc_next[7]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \input_a~144 (
// Equation(s):
// \input_a~144_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_6))) # (!MemToReg_MEM1 & (CalcData_MEM_6))))

	.dataa(\PR|CalcData_MEM [6]),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [6]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~144_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~144 .lut_mask = 16'hC088;
defparam \input_a~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \pc_next[6]~28 (
// Equation(s):
// \pc_next[6]~28_combout  = (\pc_next[6]~27_combout  & (((Result_EX_6)) # (!\pc[22]~34_combout ))) # (!\pc_next[6]~27_combout  & (\pc[22]~34_combout  & ((\input_a~144_combout ))))

	.dataa(\pc_next[6]~27_combout ),
	.datab(\pc[22]~34_combout ),
	.datac(Result_EX_6),
	.datad(\input_a~144_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~28 .lut_mask = 16'hE6A2;
defparam \pc_next[6]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \pc_next[6]~29 (
// Equation(s):
// \pc_next[6]~29_combout  = (\pc[22]~28_combout  & (\pc_next_branch[6]~8_combout )) # (!\pc[22]~28_combout  & ((\pc_next[6]~28_combout )))

	.dataa(\pc[22]~28_combout ),
	.datab(gnd),
	.datac(\pc_next_branch[6]~8_combout ),
	.datad(\pc_next[6]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~29 .lut_mask = 16'hF5A0;
defparam \pc_next[6]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \pc_next[6]~30 (
// Equation(s):
// \pc_next[6]~30_combout  = (\pc_next_plus4[6]~8_combout  & (((\pc_next[6]~29_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[6]~8_combout  & (\pc_next[6]~29_combout  & ((!\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[6]~8_combout ),
	.datab(\pc_next[6]~29_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~30 .lut_mask = 16'h0ACE;
defparam \pc_next[6]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \pc_next[9]~31 (
// Equation(s):
// \pc_next[9]~31_combout  = (\pc[22]~34_combout  & ((\input_a~145_combout ) # ((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & (((ALUSrc1_ID_9 & !\pc[22]~38_combout ))))

	.dataa(\input_a~145_combout ),
	.datab(\PR|ALUSrc1_ID [9]),
	.datac(\pc[22]~34_combout ),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~31 .lut_mask = 16'hF0AC;
defparam \pc_next[9]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \pc_next[9]~32 (
// Equation(s):
// \pc_next[9]~32_combout  = (\pc_next[9]~31_combout  & (((Result_EX_9) # (!\pc[22]~38_combout )))) # (!\pc_next[9]~31_combout  & (Instr_ID_7 & ((\pc[22]~38_combout ))))

	.dataa(\PR|Instr_ID [7]),
	.datab(\pc_next[9]~31_combout ),
	.datac(Result_EX_9),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~32_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~32 .lut_mask = 16'hE2CC;
defparam \pc_next[9]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \pc_next_branch[9]~14 (
// Equation(s):
// \pc_next_branch[9]~14_combout  = (nextPC_ID_9 & ((Instr_ID_7 & (\pc_next_branch[8]~13  & VCC)) # (!Instr_ID_7 & (!\pc_next_branch[8]~13 )))) # (!nextPC_ID_9 & ((Instr_ID_7 & (!\pc_next_branch[8]~13 )) # (!Instr_ID_7 & ((\pc_next_branch[8]~13 ) # (GND)))))
// \pc_next_branch[9]~15  = CARRY((nextPC_ID_9 & (!Instr_ID_7 & !\pc_next_branch[8]~13 )) # (!nextPC_ID_9 & ((!\pc_next_branch[8]~13 ) # (!Instr_ID_7))))

	.dataa(\PR|nextPC_ID [9]),
	.datab(\PR|Instr_ID [7]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[8]~13 ),
	.combout(\pc_next_branch[9]~14_combout ),
	.cout(\pc_next_branch[9]~15 ));
// synopsys translate_off
defparam \pc_next_branch[9]~14 .lut_mask = 16'h9617;
defparam \pc_next_branch[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \pc_next[9]~33 (
// Equation(s):
// \pc_next[9]~33_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[9]~14_combout ))) # (!\pc[22]~28_combout  & (\pc_next[9]~32_combout ))

	.dataa(gnd),
	.datab(\pc[22]~28_combout ),
	.datac(\pc_next[9]~32_combout ),
	.datad(\pc_next_branch[9]~14_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~33_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~33 .lut_mask = 16'hFC30;
defparam \pc_next[9]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \pc_next_plus4[8]~12 (
// Equation(s):
// \pc_next_plus4[8]~12_combout  = (pc_8 & (\pc_next_plus4[7]~11  $ (GND))) # (!pc_8 & (!\pc_next_plus4[7]~11  & VCC))
// \pc_next_plus4[8]~13  = CARRY((pc_8 & !\pc_next_plus4[7]~11 ))

	.dataa(pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[7]~11 ),
	.combout(\pc_next_plus4[8]~12_combout ),
	.cout(\pc_next_plus4[8]~13 ));
// synopsys translate_off
defparam \pc_next_plus4[8]~12 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \pc_next_plus4[9]~14 (
// Equation(s):
// \pc_next_plus4[9]~14_combout  = (pc_9 & (!\pc_next_plus4[8]~13 )) # (!pc_9 & ((\pc_next_plus4[8]~13 ) # (GND)))
// \pc_next_plus4[9]~15  = CARRY((!\pc_next_plus4[8]~13 ) # (!pc_9))

	.dataa(gnd),
	.datab(pc_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[8]~13 ),
	.combout(\pc_next_plus4[9]~14_combout ),
	.cout(\pc_next_plus4[9]~15 ));
// synopsys translate_off
defparam \pc_next_plus4[9]~14 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \pc_next[9]~34 (
// Equation(s):
// \pc_next[9]~34_combout  = (\pc_next[9]~33_combout  & (((!\pc[1]~26_combout  & \pc_next_plus4[9]~14_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[9]~33_combout  & (!\pc[1]~26_combout  & (\pc_next_plus4[9]~14_combout )))

	.dataa(\pc_next[9]~33_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next_plus4[9]~14_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~34_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~34 .lut_mask = 16'h30BA;
defparam \pc_next[9]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \pc_next[8]~35 (
// Equation(s):
// \pc_next[8]~35_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & (Instr_ID_6)) # (!\pc[22]~38_combout  & ((ALUSrc1_ID_8)))))

	.dataa(\PR|Instr_ID [6]),
	.datab(\pc[22]~34_combout ),
	.datac(\PR|ALUSrc1_ID [8]),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~35_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~35 .lut_mask = 16'hEE30;
defparam \pc_next[8]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \input_a~146 (
// Equation(s):
// \input_a~146_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_8)) # (!MemToReg_MEM1 & ((CalcData_MEM_8)))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|ReadData_MEM [8]),
	.datac(\PR|CalcData_MEM [8]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~146_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~146 .lut_mask = 16'h88A0;
defparam \input_a~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \pc_next[8]~36 (
// Equation(s):
// \pc_next[8]~36_combout  = (\pc[22]~34_combout  & ((\pc_next[8]~35_combout  & (Result_EX_8)) # (!\pc_next[8]~35_combout  & ((\input_a~146_combout ))))) # (!\pc[22]~34_combout  & (((\pc_next[8]~35_combout ))))

	.dataa(Result_EX_8),
	.datab(\pc[22]~34_combout ),
	.datac(\pc_next[8]~35_combout ),
	.datad(\input_a~146_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~36_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~36 .lut_mask = 16'hBCB0;
defparam \pc_next[8]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \pc_next[8]~37 (
// Equation(s):
// \pc_next[8]~37_combout  = (\pc[22]~28_combout  & (\pc_next_branch[8]~12_combout )) # (!\pc[22]~28_combout  & ((\pc_next[8]~36_combout )))

	.dataa(\pc_next_branch[8]~12_combout ),
	.datab(\pc_next[8]~36_combout ),
	.datac(gnd),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~37_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~37 .lut_mask = 16'hAACC;
defparam \pc_next[8]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \pc_next[8]~38 (
// Equation(s):
// \pc_next[8]~38_combout  = (\pc_next[8]~37_combout  & (((!\pc[1]~26_combout  & \pc_next_plus4[8]~12_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[8]~37_combout  & (!\pc[1]~26_combout  & (\pc_next_plus4[8]~12_combout )))

	.dataa(\pc_next[8]~37_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next_plus4[8]~12_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~38_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~38 .lut_mask = 16'h30BA;
defparam \pc_next[8]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N18
cycloneive_lcell_comb \pc_next_plus4[10]~16 (
// Equation(s):
// \pc_next_plus4[10]~16_combout  = (pc_10 & (\pc_next_plus4[9]~15  $ (GND))) # (!pc_10 & (!\pc_next_plus4[9]~15  & VCC))
// \pc_next_plus4[10]~17  = CARRY((pc_10 & !\pc_next_plus4[9]~15 ))

	.dataa(gnd),
	.datab(pc_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[9]~15 ),
	.combout(\pc_next_plus4[10]~16_combout ),
	.cout(\pc_next_plus4[10]~17 ));
// synopsys translate_off
defparam \pc_next_plus4[10]~16 .lut_mask = 16'hC30C;
defparam \pc_next_plus4[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \pc_next_plus4[11]~18 (
// Equation(s):
// \pc_next_plus4[11]~18_combout  = (pc_11 & (!\pc_next_plus4[10]~17 )) # (!pc_11 & ((\pc_next_plus4[10]~17 ) # (GND)))
// \pc_next_plus4[11]~19  = CARRY((!\pc_next_plus4[10]~17 ) # (!pc_11))

	.dataa(gnd),
	.datab(pc_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[10]~17 ),
	.combout(\pc_next_plus4[11]~18_combout ),
	.cout(\pc_next_plus4[11]~19 ));
// synopsys translate_off
defparam \pc_next_plus4[11]~18 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N4
cycloneive_lcell_comb \input_a~147 (
// Equation(s):
// \input_a~147_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_11)) # (!MemToReg_MEM1 & ((CalcData_MEM_11)))))

	.dataa(\PR|ReadData_MEM [11]),
	.datab(\PR|CalcData_MEM [11]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~147_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~147 .lut_mask = 16'hA0C0;
defparam \input_a~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \pc_next[11]~39 (
// Equation(s):
// \pc_next[11]~39_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & ((\input_a~147_combout ))) # (!\pc[22]~34_combout  & (ALUSrc1_ID_11))))

	.dataa(\PR|ALUSrc1_ID [11]),
	.datab(\input_a~147_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~39_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~39 .lut_mask = 16'hFC0A;
defparam \pc_next[11]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \pc_next[11]~40 (
// Equation(s):
// \pc_next[11]~40_combout  = (\pc[22]~38_combout  & ((\pc_next[11]~39_combout  & (Result_EX_11)) # (!\pc_next[11]~39_combout  & ((Instr_ID_9))))) # (!\pc[22]~38_combout  & (((\pc_next[11]~39_combout ))))

	.dataa(Result_EX_11),
	.datab(\PR|Instr_ID [9]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc_next[11]~39_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~40_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~40 .lut_mask = 16'hAFC0;
defparam \pc_next[11]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \pc_next_branch[10]~16 (
// Equation(s):
// \pc_next_branch[10]~16_combout  = ((Instr_ID_8 $ (nextPC_ID_10 $ (!\pc_next_branch[9]~15 )))) # (GND)
// \pc_next_branch[10]~17  = CARRY((Instr_ID_8 & ((nextPC_ID_10) # (!\pc_next_branch[9]~15 ))) # (!Instr_ID_8 & (nextPC_ID_10 & !\pc_next_branch[9]~15 )))

	.dataa(\PR|Instr_ID [8]),
	.datab(\PR|nextPC_ID [10]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[9]~15 ),
	.combout(\pc_next_branch[10]~16_combout ),
	.cout(\pc_next_branch[10]~17 ));
// synopsys translate_off
defparam \pc_next_branch[10]~16 .lut_mask = 16'h698E;
defparam \pc_next_branch[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \pc_next_branch[11]~18 (
// Equation(s):
// \pc_next_branch[11]~18_combout  = (Instr_ID_9 & ((nextPC_ID_11 & (\pc_next_branch[10]~17  & VCC)) # (!nextPC_ID_11 & (!\pc_next_branch[10]~17 )))) # (!Instr_ID_9 & ((nextPC_ID_11 & (!\pc_next_branch[10]~17 )) # (!nextPC_ID_11 & ((\pc_next_branch[10]~17 ) 
// # (GND)))))
// \pc_next_branch[11]~19  = CARRY((Instr_ID_9 & (!nextPC_ID_11 & !\pc_next_branch[10]~17 )) # (!Instr_ID_9 & ((!\pc_next_branch[10]~17 ) # (!nextPC_ID_11))))

	.dataa(\PR|Instr_ID [9]),
	.datab(\PR|nextPC_ID [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[10]~17 ),
	.combout(\pc_next_branch[11]~18_combout ),
	.cout(\pc_next_branch[11]~19 ));
// synopsys translate_off
defparam \pc_next_branch[11]~18 .lut_mask = 16'h9617;
defparam \pc_next_branch[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \pc_next[11]~41 (
// Equation(s):
// \pc_next[11]~41_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[11]~18_combout ))) # (!\pc[22]~28_combout  & (\pc_next[11]~40_combout ))

	.dataa(\pc[22]~28_combout ),
	.datab(gnd),
	.datac(\pc_next[11]~40_combout ),
	.datad(\pc_next_branch[11]~18_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~41_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~41 .lut_mask = 16'hFA50;
defparam \pc_next[11]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \pc_next[11]~42 (
// Equation(s):
// \pc_next[11]~42_combout  = (\pc_next_plus4[11]~18_combout  & (((\pc_next[11]~41_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[11]~18_combout  & (((\pc_next[11]~41_combout  & !\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[11]~18_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next[11]~41_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~42_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~42 .lut_mask = 16'h22F2;
defparam \pc_next[11]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \pc_next[10]~43 (
// Equation(s):
// \pc_next[10]~43_combout  = (\pc[22]~38_combout  & ((Instr_ID_8) # ((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (((ALUSrc1_ID_10 & !\pc[22]~34_combout ))))

	.dataa(\PR|Instr_ID [8]),
	.datab(\PR|ALUSrc1_ID [10]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~43_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~43 .lut_mask = 16'hF0AC;
defparam \pc_next[10]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N30
cycloneive_lcell_comb \input_a~148 (
// Equation(s):
// \input_a~148_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_10))) # (!MemToReg_MEM1 & (CalcData_MEM_10))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|CalcData_MEM [10]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|ReadData_MEM [10]),
	.cin(gnd),
	.combout(\input_a~148_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~148 .lut_mask = 16'hA808;
defparam \input_a~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \pc_next[10]~44 (
// Equation(s):
// \pc_next[10]~44_combout  = (\pc[22]~34_combout  & ((\pc_next[10]~43_combout  & (Result_EX_10)) # (!\pc_next[10]~43_combout  & ((\input_a~148_combout ))))) # (!\pc[22]~34_combout  & (\pc_next[10]~43_combout ))

	.dataa(\pc[22]~34_combout ),
	.datab(\pc_next[10]~43_combout ),
	.datac(Result_EX_10),
	.datad(\input_a~148_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~44_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~44 .lut_mask = 16'hE6C4;
defparam \pc_next[10]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \pc_next[10]~45 (
// Equation(s):
// \pc_next[10]~45_combout  = (\pc[22]~28_combout  & (\pc_next_branch[10]~16_combout )) # (!\pc[22]~28_combout  & ((\pc_next[10]~44_combout )))

	.dataa(\pc[22]~28_combout ),
	.datab(\pc_next_branch[10]~16_combout ),
	.datac(\pc_next[10]~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_next[10]~45_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~45 .lut_mask = 16'hD8D8;
defparam \pc_next[10]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \pc_next[10]~46 (
// Equation(s):
// \pc_next[10]~46_combout  = (\pc_next_plus4[10]~16_combout  & (((\pc_next[10]~45_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[10]~16_combout  & (\pc_next[10]~45_combout  & ((!\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[10]~16_combout ),
	.datab(\pc_next[10]~45_combout ),
	.datac(\pc[1]~26_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~46_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~46 .lut_mask = 16'h0ACE;
defparam \pc_next[10]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \pc_next_plus4[12]~20 (
// Equation(s):
// \pc_next_plus4[12]~20_combout  = (pc_12 & (\pc_next_plus4[11]~19  $ (GND))) # (!pc_12 & (!\pc_next_plus4[11]~19  & VCC))
// \pc_next_plus4[12]~21  = CARRY((pc_12 & !\pc_next_plus4[11]~19 ))

	.dataa(gnd),
	.datab(pc_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[11]~19 ),
	.combout(\pc_next_plus4[12]~20_combout ),
	.cout(\pc_next_plus4[12]~21 ));
// synopsys translate_off
defparam \pc_next_plus4[12]~20 .lut_mask = 16'hC30C;
defparam \pc_next_plus4[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \pc_next_plus4[13]~22 (
// Equation(s):
// \pc_next_plus4[13]~22_combout  = (pc_13 & (!\pc_next_plus4[12]~21 )) # (!pc_13 & ((\pc_next_plus4[12]~21 ) # (GND)))
// \pc_next_plus4[13]~23  = CARRY((!\pc_next_plus4[12]~21 ) # (!pc_13))

	.dataa(gnd),
	.datab(pc_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[12]~21 ),
	.combout(\pc_next_plus4[13]~22_combout ),
	.cout(\pc_next_plus4[13]~23 ));
// synopsys translate_off
defparam \pc_next_plus4[13]~22 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \pc_next_branch[12]~20 (
// Equation(s):
// \pc_next_branch[12]~20_combout  = ((Instr_ID_10 $ (nextPC_ID_12 $ (!\pc_next_branch[11]~19 )))) # (GND)
// \pc_next_branch[12]~21  = CARRY((Instr_ID_10 & ((nextPC_ID_12) # (!\pc_next_branch[11]~19 ))) # (!Instr_ID_10 & (nextPC_ID_12 & !\pc_next_branch[11]~19 )))

	.dataa(\PR|Instr_ID [10]),
	.datab(\PR|nextPC_ID [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[11]~19 ),
	.combout(\pc_next_branch[12]~20_combout ),
	.cout(\pc_next_branch[12]~21 ));
// synopsys translate_off
defparam \pc_next_branch[12]~20 .lut_mask = 16'h698E;
defparam \pc_next_branch[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \pc_next_branch[13]~22 (
// Equation(s):
// \pc_next_branch[13]~22_combout  = (nextPC_ID_13 & ((Instr_ID_11 & (\pc_next_branch[12]~21  & VCC)) # (!Instr_ID_11 & (!\pc_next_branch[12]~21 )))) # (!nextPC_ID_13 & ((Instr_ID_11 & (!\pc_next_branch[12]~21 )) # (!Instr_ID_11 & ((\pc_next_branch[12]~21 ) 
// # (GND)))))
// \pc_next_branch[13]~23  = CARRY((nextPC_ID_13 & (!Instr_ID_11 & !\pc_next_branch[12]~21 )) # (!nextPC_ID_13 & ((!\pc_next_branch[12]~21 ) # (!Instr_ID_11))))

	.dataa(\PR|nextPC_ID [13]),
	.datab(\PR|Instr_ID [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[12]~21 ),
	.combout(\pc_next_branch[13]~22_combout ),
	.cout(\pc_next_branch[13]~23 ));
// synopsys translate_off
defparam \pc_next_branch[13]~22 .lut_mask = 16'h9617;
defparam \pc_next_branch[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \input_a~149 (
// Equation(s):
// \input_a~149_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_13)) # (!MemToReg_MEM1 & ((CalcData_MEM_13)))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|ReadData_MEM [13]),
	.datac(\PR|CalcData_MEM [13]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~149_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~149 .lut_mask = 16'h88A0;
defparam \input_a~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \pc_next[13]~47 (
// Equation(s):
// \pc_next[13]~47_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & (\input_a~149_combout )) # (!\pc[22]~34_combout  & ((ALUSrc1_ID_13)))))

	.dataa(\pc[22]~38_combout ),
	.datab(\input_a~149_combout ),
	.datac(\PR|ALUSrc1_ID [13]),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~47_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~47 .lut_mask = 16'hEE50;
defparam \pc_next[13]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \pc_next[13]~48 (
// Equation(s):
// \pc_next[13]~48_combout  = (\pc[22]~38_combout  & ((\pc_next[13]~47_combout  & ((Result_EX_13))) # (!\pc_next[13]~47_combout  & (Instr_ID_11)))) # (!\pc[22]~38_combout  & (((\pc_next[13]~47_combout ))))

	.dataa(\pc[22]~38_combout ),
	.datab(\PR|Instr_ID [11]),
	.datac(Result_EX_13),
	.datad(\pc_next[13]~47_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~48_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~48 .lut_mask = 16'hF588;
defparam \pc_next[13]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N4
cycloneive_lcell_comb \pc_next[13]~49 (
// Equation(s):
// \pc_next[13]~49_combout  = (\pc[22]~28_combout  & (\pc_next_branch[13]~22_combout )) # (!\pc[22]~28_combout  & ((\pc_next[13]~48_combout )))

	.dataa(gnd),
	.datab(\pc[22]~28_combout ),
	.datac(\pc_next_branch[13]~22_combout ),
	.datad(\pc_next[13]~48_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~49_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~49 .lut_mask = 16'hF3C0;
defparam \pc_next[13]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N8
cycloneive_lcell_comb \pc_next[13]~50 (
// Equation(s):
// \pc_next[13]~50_combout  = (\pc_next_plus4[13]~22_combout  & (((\pc_next[13]~49_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[13]~22_combout  & (((\pc_next[13]~49_combout  & !\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[13]~22_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next[13]~49_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~50_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~50 .lut_mask = 16'h22F2;
defparam \pc_next[13]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N28
cycloneive_lcell_comb \input_a~150 (
// Equation(s):
// \input_a~150_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_12))) # (!MemToReg_MEM1 & (CalcData_MEM_12))))

	.dataa(\PR|CalcData_MEM [12]),
	.datab(\PR|MemToReg_MEM~q ),
	.datac(\PR|ReadData_MEM [12]),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~150_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~150 .lut_mask = 16'hE200;
defparam \input_a~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \pc_next[12]~51 (
// Equation(s):
// \pc_next[12]~51_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & (Instr_ID_10)) # (!\pc[22]~38_combout  & ((ALUSrc1_ID_12)))))

	.dataa(\pc[22]~34_combout ),
	.datab(\PR|Instr_ID [10]),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|ALUSrc1_ID [12]),
	.cin(gnd),
	.combout(\pc_next[12]~51_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~51 .lut_mask = 16'hE5E0;
defparam \pc_next[12]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N8
cycloneive_lcell_comb \pc_next[12]~52 (
// Equation(s):
// \pc_next[12]~52_combout  = (\pc_next[12]~51_combout  & ((Result_EX_12) # ((!\pc[22]~34_combout )))) # (!\pc_next[12]~51_combout  & (((\input_a~150_combout  & \pc[22]~34_combout ))))

	.dataa(Result_EX_12),
	.datab(\input_a~150_combout ),
	.datac(\pc_next[12]~51_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[12]~52_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~52 .lut_mask = 16'hACF0;
defparam \pc_next[12]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N2
cycloneive_lcell_comb \pc_next[12]~53 (
// Equation(s):
// \pc_next[12]~53_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[12]~20_combout ))) # (!\pc[22]~28_combout  & (\pc_next[12]~52_combout ))

	.dataa(gnd),
	.datab(\pc_next[12]~52_combout ),
	.datac(\pc[22]~28_combout ),
	.datad(\pc_next_branch[12]~20_combout ),
	.cin(gnd),
	.combout(\pc_next[12]~53_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~53 .lut_mask = 16'hFC0C;
defparam \pc_next[12]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N4
cycloneive_lcell_comb \pc_next[12]~54 (
// Equation(s):
// \pc_next[12]~54_combout  = (\pc_next[12]~53_combout  & (((!\pc[1]~26_combout  & \pc_next_plus4[12]~20_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[12]~53_combout  & (!\pc[1]~26_combout  & (\pc_next_plus4[12]~20_combout )))

	.dataa(\pc_next[12]~53_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next_plus4[12]~20_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[12]~54_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~54 .lut_mask = 16'h30BA;
defparam \pc_next[12]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \input_a~151 (
// Equation(s):
// \input_a~151_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_15)) # (!MemToReg_MEM1 & ((CalcData_MEM_15)))))

	.dataa(\PR|ReadData_MEM [15]),
	.datab(\PR|CalcData_MEM [15]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~151_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~151 .lut_mask = 16'hA0C0;
defparam \input_a~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N6
cycloneive_lcell_comb \pc_next[15]~55 (
// Equation(s):
// \pc_next[15]~55_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & ((\input_a~151_combout ))) # (!\pc[22]~34_combout  & (ALUSrc1_ID_15))))

	.dataa(\PR|ALUSrc1_ID [15]),
	.datab(\input_a~151_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~55_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~55 .lut_mask = 16'hFC0A;
defparam \pc_next[15]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N16
cycloneive_lcell_comb \pc_next[15]~56 (
// Equation(s):
// \pc_next[15]~56_combout  = (\pc_next[15]~55_combout  & ((Result_EX_15) # ((!\pc[22]~38_combout )))) # (!\pc_next[15]~55_combout  & (((Instr_ID_13 & \pc[22]~38_combout ))))

	.dataa(Result_EX_15),
	.datab(\PR|Instr_ID [13]),
	.datac(\pc_next[15]~55_combout ),
	.datad(\pc[22]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~56_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~56 .lut_mask = 16'hACF0;
defparam \pc_next[15]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \pc_next_branch[14]~24 (
// Equation(s):
// \pc_next_branch[14]~24_combout  = ((nextPC_ID_14 $ (Instr_ID_12 $ (!\pc_next_branch[13]~23 )))) # (GND)
// \pc_next_branch[14]~25  = CARRY((nextPC_ID_14 & ((Instr_ID_12) # (!\pc_next_branch[13]~23 ))) # (!nextPC_ID_14 & (Instr_ID_12 & !\pc_next_branch[13]~23 )))

	.dataa(\PR|nextPC_ID [14]),
	.datab(\PR|Instr_ID [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[13]~23 ),
	.combout(\pc_next_branch[14]~24_combout ),
	.cout(\pc_next_branch[14]~25 ));
// synopsys translate_off
defparam \pc_next_branch[14]~24 .lut_mask = 16'h698E;
defparam \pc_next_branch[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \pc_next_branch[15]~26 (
// Equation(s):
// \pc_next_branch[15]~26_combout  = (Instr_ID_13 & ((nextPC_ID_15 & (\pc_next_branch[14]~25  & VCC)) # (!nextPC_ID_15 & (!\pc_next_branch[14]~25 )))) # (!Instr_ID_13 & ((nextPC_ID_15 & (!\pc_next_branch[14]~25 )) # (!nextPC_ID_15 & ((\pc_next_branch[14]~25 
// ) # (GND)))))
// \pc_next_branch[15]~27  = CARRY((Instr_ID_13 & (!nextPC_ID_15 & !\pc_next_branch[14]~25 )) # (!Instr_ID_13 & ((!\pc_next_branch[14]~25 ) # (!nextPC_ID_15))))

	.dataa(\PR|Instr_ID [13]),
	.datab(\PR|nextPC_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[14]~25 ),
	.combout(\pc_next_branch[15]~26_combout ),
	.cout(\pc_next_branch[15]~27 ));
// synopsys translate_off
defparam \pc_next_branch[15]~26 .lut_mask = 16'h9617;
defparam \pc_next_branch[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N2
cycloneive_lcell_comb \pc_next[15]~57 (
// Equation(s):
// \pc_next[15]~57_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[15]~26_combout ))) # (!\pc[22]~28_combout  & (\pc_next[15]~56_combout ))

	.dataa(gnd),
	.datab(\pc_next[15]~56_combout ),
	.datac(\pc_next_branch[15]~26_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~57_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~57 .lut_mask = 16'hF0CC;
defparam \pc_next[15]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \pc_next_plus4[14]~24 (
// Equation(s):
// \pc_next_plus4[14]~24_combout  = (pc_14 & (\pc_next_plus4[13]~23  $ (GND))) # (!pc_14 & (!\pc_next_plus4[13]~23  & VCC))
// \pc_next_plus4[14]~25  = CARRY((pc_14 & !\pc_next_plus4[13]~23 ))

	.dataa(pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[13]~23 ),
	.combout(\pc_next_plus4[14]~24_combout ),
	.cout(\pc_next_plus4[14]~25 ));
// synopsys translate_off
defparam \pc_next_plus4[14]~24 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \pc_next_plus4[15]~26 (
// Equation(s):
// \pc_next_plus4[15]~26_combout  = (pc_15 & (!\pc_next_plus4[14]~25 )) # (!pc_15 & ((\pc_next_plus4[14]~25 ) # (GND)))
// \pc_next_plus4[15]~27  = CARRY((!\pc_next_plus4[14]~25 ) # (!pc_15))

	.dataa(pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[14]~25 ),
	.combout(\pc_next_plus4[15]~26_combout ),
	.cout(\pc_next_plus4[15]~27 ));
// synopsys translate_off
defparam \pc_next_plus4[15]~26 .lut_mask = 16'h5A5F;
defparam \pc_next_plus4[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N8
cycloneive_lcell_comb \pc_next[15]~58 (
// Equation(s):
// \pc_next[15]~58_combout  = (\pc_next[15]~57_combout  & (((\pc_next_plus4[15]~26_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[15]~57_combout  & (\pc_next_plus4[15]~26_combout  & ((!\pc[1]~26_combout ))))

	.dataa(\pc_next[15]~57_combout ),
	.datab(\pc_next_plus4[15]~26_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~58 .lut_mask = 16'h0ACE;
defparam \pc_next[15]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N14
cycloneive_lcell_comb \pc_next[14]~59 (
// Equation(s):
// \pc_next[14]~59_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & (Instr_ID_12)) # (!\pc[22]~38_combout  & ((ALUSrc1_ID_14)))))

	.dataa(\pc[22]~34_combout ),
	.datab(\PR|Instr_ID [12]),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|ALUSrc1_ID [14]),
	.cin(gnd),
	.combout(\pc_next[14]~59_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~59 .lut_mask = 16'hE5E0;
defparam \pc_next[14]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \pc_next[14]~60 (
// Equation(s):
// \pc_next[14]~60_combout  = (\pc_next[14]~59_combout  & (((Result_EX_14) # (!\pc[22]~34_combout )))) # (!\pc_next[14]~59_combout  & (\input_a~152_combout  & ((\pc[22]~34_combout ))))

	.dataa(\input_a~152_combout ),
	.datab(\pc_next[14]~59_combout ),
	.datac(Result_EX_14),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[14]~60_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~60 .lut_mask = 16'hE2CC;
defparam \pc_next[14]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N20
cycloneive_lcell_comb \pc_next[14]~61 (
// Equation(s):
// \pc_next[14]~61_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[14]~24_combout ))) # (!\pc[22]~28_combout  & (\pc_next[14]~60_combout ))

	.dataa(\pc[22]~28_combout ),
	.datab(gnd),
	.datac(\pc_next[14]~60_combout ),
	.datad(\pc_next_branch[14]~24_combout ),
	.cin(gnd),
	.combout(\pc_next[14]~61_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~61 .lut_mask = 16'hFA50;
defparam \pc_next[14]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \pc_next[14]~62 (
// Equation(s):
// \pc_next[14]~62_combout  = (\pc_next_plus4[14]~24_combout  & (((\pc_next[14]~61_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[14]~24_combout  & (((\pc_next[14]~61_combout  & !\pc_next[27]~9_combout ))))

	.dataa(\pc_next_plus4[14]~24_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next[14]~61_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[14]~62_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~62 .lut_mask = 16'h22F2;
defparam \pc_next[14]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \pc_next_plus4[16]~28 (
// Equation(s):
// \pc_next_plus4[16]~28_combout  = (pc_16 & (\pc_next_plus4[15]~27  $ (GND))) # (!pc_16 & (!\pc_next_plus4[15]~27  & VCC))
// \pc_next_plus4[16]~29  = CARRY((pc_16 & !\pc_next_plus4[15]~27 ))

	.dataa(gnd),
	.datab(pc_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[15]~27 ),
	.combout(\pc_next_plus4[16]~28_combout ),
	.cout(\pc_next_plus4[16]~29 ));
// synopsys translate_off
defparam \pc_next_plus4[16]~28 .lut_mask = 16'hC30C;
defparam \pc_next_plus4[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N0
cycloneive_lcell_comb \pc_next_plus4[17]~30 (
// Equation(s):
// \pc_next_plus4[17]~30_combout  = (pc_17 & (!\pc_next_plus4[16]~29 )) # (!pc_17 & ((\pc_next_plus4[16]~29 ) # (GND)))
// \pc_next_plus4[17]~31  = CARRY((!\pc_next_plus4[16]~29 ) # (!pc_17))

	.dataa(gnd),
	.datab(pc_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[16]~29 ),
	.combout(\pc_next_plus4[17]~30_combout ),
	.cout(\pc_next_plus4[17]~31 ));
// synopsys translate_off
defparam \pc_next_plus4[17]~30 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \input_a~153 (
// Equation(s):
// \input_a~153_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_17))) # (!MemToReg_MEM1 & (CalcData_MEM_17))))

	.dataa(\PR|CalcData_MEM [17]),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [17]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~153_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~153 .lut_mask = 16'hC088;
defparam \input_a~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \pc_next[17]~63 (
// Equation(s):
// \pc_next[17]~63_combout  = (\pc[22]~34_combout  & ((\pc[22]~38_combout ) # ((\input_a~153_combout )))) # (!\pc[22]~34_combout  & (!\pc[22]~38_combout  & ((ALUSrc1_ID_17))))

	.dataa(\pc[22]~34_combout ),
	.datab(\pc[22]~38_combout ),
	.datac(\input_a~153_combout ),
	.datad(\PR|ALUSrc1_ID [17]),
	.cin(gnd),
	.combout(\pc_next[17]~63_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~63 .lut_mask = 16'hB9A8;
defparam \pc_next[17]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \pc_next[17]~64 (
// Equation(s):
// \pc_next[17]~64_combout  = (\pc[22]~38_combout  & ((\pc_next[17]~63_combout  & ((Result_EX_17))) # (!\pc_next[17]~63_combout  & (Instr_ID_15)))) # (!\pc[22]~38_combout  & (((\pc_next[17]~63_combout ))))

	.dataa(\PR|Instr_ID [15]),
	.datab(\pc[22]~38_combout ),
	.datac(Result_EX_17),
	.datad(\pc_next[17]~63_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~64_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~64 .lut_mask = 16'hF388;
defparam \pc_next[17]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \pc_next[17]~65 (
// Equation(s):
// \pc_next[17]~65_combout  = (\pc[22]~28_combout  & (\pc_next_branch[17]~30_combout )) # (!\pc[22]~28_combout  & ((\pc_next[17]~64_combout )))

	.dataa(\pc_next_branch[17]~30_combout ),
	.datab(\pc_next[17]~64_combout ),
	.datac(gnd),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~65_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~65 .lut_mask = 16'hAACC;
defparam \pc_next[17]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \pc_next[17]~66 (
// Equation(s):
// \pc_next[17]~66_combout  = (\pc_next_plus4[17]~30_combout  & (((\pc_next[17]~65_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[17]~30_combout  & (\pc_next[17]~65_combout  & (!\pc_next[27]~9_combout )))

	.dataa(\pc_next_plus4[17]~30_combout ),
	.datab(\pc_next[17]~65_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~66_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~66 .lut_mask = 16'h0CAE;
defparam \pc_next[17]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \input_a~154 (
// Equation(s):
// \input_a~154_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_16)) # (!MemToReg_MEM1 & ((CalcData_MEM_16)))))

	.dataa(\Equal24~0_combout ),
	.datab(\PR|ReadData_MEM [16]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\PR|CalcData_MEM [16]),
	.cin(gnd),
	.combout(\input_a~154_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~154 .lut_mask = 16'h8A80;
defparam \input_a~154 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \pc_next[16]~67 (
// Equation(s):
// \pc_next[16]~67_combout  = (\pc[22]~38_combout  & ((Instr_ID_14) # ((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (((ALUSrc1_ID_16 & !\pc[22]~34_combout ))))

	.dataa(\PR|Instr_ID [14]),
	.datab(\PR|ALUSrc1_ID [16]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~67_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~67 .lut_mask = 16'hF0AC;
defparam \pc_next[16]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \pc_next[16]~68 (
// Equation(s):
// \pc_next[16]~68_combout  = (\pc[22]~34_combout  & ((\pc_next[16]~67_combout  & ((Result_EX_16))) # (!\pc_next[16]~67_combout  & (\input_a~154_combout )))) # (!\pc[22]~34_combout  & (((\pc_next[16]~67_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(\input_a~154_combout ),
	.datac(Result_EX_16),
	.datad(\pc_next[16]~67_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~68_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~68 .lut_mask = 16'hF588;
defparam \pc_next[16]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \pc_next[16]~69 (
// Equation(s):
// \pc_next[16]~69_combout  = (\pc[22]~28_combout  & (\pc_next_branch[16]~28_combout )) # (!\pc[22]~28_combout  & ((\pc_next[16]~68_combout )))

	.dataa(\pc_next_branch[16]~28_combout ),
	.datab(\pc_next[16]~68_combout ),
	.datac(gnd),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~69_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~69 .lut_mask = 16'hAACC;
defparam \pc_next[16]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \pc_next[16]~70 (
// Equation(s):
// \pc_next[16]~70_combout  = (\pc_next_plus4[16]~28_combout  & (((\pc_next[16]~69_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[16]~28_combout  & (\pc_next[16]~69_combout  & (!\pc_next[27]~9_combout )))

	.dataa(\pc_next_plus4[16]~28_combout ),
	.datab(\pc_next[16]~69_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~70_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~70 .lut_mask = 16'h0CAE;
defparam \pc_next[16]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N4
cycloneive_lcell_comb \pc_next_branch[19]~34 (
// Equation(s):
// \pc_next_branch[19]~34_combout  = (nextPC_ID_19 & ((Instr_ID_15 & (\pc_next_branch[18]~33  & VCC)) # (!Instr_ID_15 & (!\pc_next_branch[18]~33 )))) # (!nextPC_ID_19 & ((Instr_ID_15 & (!\pc_next_branch[18]~33 )) # (!Instr_ID_15 & ((\pc_next_branch[18]~33 ) 
// # (GND)))))
// \pc_next_branch[19]~35  = CARRY((nextPC_ID_19 & (!Instr_ID_15 & !\pc_next_branch[18]~33 )) # (!nextPC_ID_19 & ((!\pc_next_branch[18]~33 ) # (!Instr_ID_15))))

	.dataa(\PR|nextPC_ID [19]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[18]~33 ),
	.combout(\pc_next_branch[19]~34_combout ),
	.cout(\pc_next_branch[19]~35 ));
// synopsys translate_off
defparam \pc_next_branch[19]~34 .lut_mask = 16'h9617;
defparam \pc_next_branch[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \pc_next[19]~73 (
// Equation(s):
// \pc_next[19]~73_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[19]~34_combout ))) # (!\pc[22]~28_combout  & (\pc_next[19]~72_combout ))

	.dataa(\pc_next[19]~72_combout ),
	.datab(gnd),
	.datac(\pc_next_branch[19]~34_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[19]~73_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~73 .lut_mask = 16'hF0AA;
defparam \pc_next[19]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N2
cycloneive_lcell_comb \pc_next_plus4[18]~32 (
// Equation(s):
// \pc_next_plus4[18]~32_combout  = (pc_18 & (\pc_next_plus4[17]~31  $ (GND))) # (!pc_18 & (!\pc_next_plus4[17]~31  & VCC))
// \pc_next_plus4[18]~33  = CARRY((pc_18 & !\pc_next_plus4[17]~31 ))

	.dataa(pc_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[17]~31 ),
	.combout(\pc_next_plus4[18]~32_combout ),
	.cout(\pc_next_plus4[18]~33 ));
// synopsys translate_off
defparam \pc_next_plus4[18]~32 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N4
cycloneive_lcell_comb \pc_next_plus4[19]~34 (
// Equation(s):
// \pc_next_plus4[19]~34_combout  = (pc_19 & (!\pc_next_plus4[18]~33 )) # (!pc_19 & ((\pc_next_plus4[18]~33 ) # (GND)))
// \pc_next_plus4[19]~35  = CARRY((!\pc_next_plus4[18]~33 ) # (!pc_19))

	.dataa(gnd),
	.datab(pc_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[18]~33 ),
	.combout(\pc_next_plus4[19]~34_combout ),
	.cout(\pc_next_plus4[19]~35 ));
// synopsys translate_off
defparam \pc_next_plus4[19]~34 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \pc_next[19]~74 (
// Equation(s):
// \pc_next[19]~74_combout  = (\pc[1]~26_combout  & (\pc_next[19]~73_combout  & (!\pc_next[27]~9_combout ))) # (!\pc[1]~26_combout  & ((\pc_next_plus4[19]~34_combout ) # ((\pc_next[19]~73_combout  & !\pc_next[27]~9_combout ))))

	.dataa(\pc[1]~26_combout ),
	.datab(\pc_next[19]~73_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc_next_plus4[19]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[19]~74_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~74 .lut_mask = 16'h5D0C;
defparam \pc_next[19]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \pc_next[18]~75 (
// Equation(s):
// \pc_next[18]~75_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & (Instr_ID_16)) # (!\pc[22]~38_combout  & ((ALUSrc1_ID_18)))))

	.dataa(\pc[22]~34_combout ),
	.datab(\PR|Instr_ID [16]),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|ALUSrc1_ID [18]),
	.cin(gnd),
	.combout(\pc_next[18]~75_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~75 .lut_mask = 16'hE5E0;
defparam \pc_next[18]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \input_a~156 (
// Equation(s):
// \input_a~156_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_18)) # (!MemToReg_MEM1 & ((CalcData_MEM_18)))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|ReadData_MEM [18]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|CalcData_MEM [18]),
	.cin(gnd),
	.combout(\input_a~156_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~156 .lut_mask = 16'hD080;
defparam \input_a~156 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \pc_next[18]~76 (
// Equation(s):
// \pc_next[18]~76_combout  = (\pc[22]~34_combout  & ((\pc_next[18]~75_combout  & (Result_EX_18)) # (!\pc_next[18]~75_combout  & ((\input_a~156_combout ))))) # (!\pc[22]~34_combout  & (((\pc_next[18]~75_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(Result_EX_18),
	.datac(\pc_next[18]~75_combout ),
	.datad(\input_a~156_combout ),
	.cin(gnd),
	.combout(\pc_next[18]~76_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~76 .lut_mask = 16'hDAD0;
defparam \pc_next[18]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \pc_next[18]~77 (
// Equation(s):
// \pc_next[18]~77_combout  = (\pc[22]~28_combout  & (\pc_next_branch[18]~32_combout )) # (!\pc[22]~28_combout  & ((\pc_next[18]~76_combout )))

	.dataa(\pc_next_branch[18]~32_combout ),
	.datab(\pc[22]~28_combout ),
	.datac(gnd),
	.datad(\pc_next[18]~76_combout ),
	.cin(gnd),
	.combout(\pc_next[18]~77_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~77 .lut_mask = 16'hBB88;
defparam \pc_next[18]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \pc_next[18]~78 (
// Equation(s):
// \pc_next[18]~78_combout  = (\pc_next_plus4[18]~32_combout  & (((\pc_next[18]~77_combout  & !\pc_next[27]~9_combout )) # (!\pc[1]~26_combout ))) # (!\pc_next_plus4[18]~32_combout  & (\pc_next[18]~77_combout  & (!\pc_next[27]~9_combout )))

	.dataa(\pc_next_plus4[18]~32_combout ),
	.datab(\pc_next[18]~77_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[18]~78_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~78 .lut_mask = 16'h0CAE;
defparam \pc_next[18]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N8
cycloneive_lcell_comb \pc_next_branch[21]~38 (
// Equation(s):
// \pc_next_branch[21]~38_combout  = (nextPC_ID_21 & ((Instr_ID_15 & (\pc_next_branch[20]~37  & VCC)) # (!Instr_ID_15 & (!\pc_next_branch[20]~37 )))) # (!nextPC_ID_21 & ((Instr_ID_15 & (!\pc_next_branch[20]~37 )) # (!Instr_ID_15 & ((\pc_next_branch[20]~37 ) 
// # (GND)))))
// \pc_next_branch[21]~39  = CARRY((nextPC_ID_21 & (!Instr_ID_15 & !\pc_next_branch[20]~37 )) # (!nextPC_ID_21 & ((!\pc_next_branch[20]~37 ) # (!Instr_ID_15))))

	.dataa(\PR|nextPC_ID [21]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[20]~37 ),
	.combout(\pc_next_branch[21]~38_combout ),
	.cout(\pc_next_branch[21]~39 ));
// synopsys translate_off
defparam \pc_next_branch[21]~38 .lut_mask = 16'h9617;
defparam \pc_next_branch[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N8
cycloneive_lcell_comb \pc_next[21]~81 (
// Equation(s):
// \pc_next[21]~81_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[21]~38_combout ))) # (!\pc[22]~28_combout  & (\pc_next[21]~80_combout ))

	.dataa(\pc_next[21]~80_combout ),
	.datab(\pc_next_branch[21]~38_combout ),
	.datac(gnd),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[21]~81_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~81 .lut_mask = 16'hCCAA;
defparam \pc_next[21]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N6
cycloneive_lcell_comb \pc_next_plus4[20]~36 (
// Equation(s):
// \pc_next_plus4[20]~36_combout  = (pc_20 & (\pc_next_plus4[19]~35  $ (GND))) # (!pc_20 & (!\pc_next_plus4[19]~35  & VCC))
// \pc_next_plus4[20]~37  = CARRY((pc_20 & !\pc_next_plus4[19]~35 ))

	.dataa(pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[19]~35 ),
	.combout(\pc_next_plus4[20]~36_combout ),
	.cout(\pc_next_plus4[20]~37 ));
// synopsys translate_off
defparam \pc_next_plus4[20]~36 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N8
cycloneive_lcell_comb \pc_next_plus4[21]~38 (
// Equation(s):
// \pc_next_plus4[21]~38_combout  = (pc_21 & (!\pc_next_plus4[20]~37 )) # (!pc_21 & ((\pc_next_plus4[20]~37 ) # (GND)))
// \pc_next_plus4[21]~39  = CARRY((!\pc_next_plus4[20]~37 ) # (!pc_21))

	.dataa(gnd),
	.datab(pc_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[20]~37 ),
	.combout(\pc_next_plus4[21]~38_combout ),
	.cout(\pc_next_plus4[21]~39 ));
// synopsys translate_off
defparam \pc_next_plus4[21]~38 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N20
cycloneive_lcell_comb \pc_next[21]~82 (
// Equation(s):
// \pc_next[21]~82_combout  = (\pc_next[21]~81_combout  & (((\pc_next_plus4[21]~38_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[21]~81_combout  & (((\pc_next_plus4[21]~38_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[21]~81_combout ),
	.datab(\pc_next[27]~9_combout ),
	.datac(\pc_next_plus4[21]~38_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[21]~82_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~82 .lut_mask = 16'h22F2;
defparam \pc_next[21]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \pc_next[20]~83 (
// Equation(s):
// \pc_next[20]~83_combout  = (\pc[22]~34_combout  & (\pc[22]~38_combout )) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & ((Instr_ID_18))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_20))))

	.dataa(\pc[22]~34_combout ),
	.datab(\pc[22]~38_combout ),
	.datac(\PR|ALUSrc1_ID [20]),
	.datad(\PR|Instr_ID [18]),
	.cin(gnd),
	.combout(\pc_next[20]~83_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~83 .lut_mask = 16'hDC98;
defparam \pc_next[20]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \input_a~158 (
// Equation(s):
// \input_a~158_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_20))) # (!MemToReg_MEM1 & (CalcData_MEM_20))))

	.dataa(\PR|CalcData_MEM [20]),
	.datab(\PR|ReadData_MEM [20]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~158_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~158 .lut_mask = 16'hC0A0;
defparam \input_a~158 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \pc_next[20]~84 (
// Equation(s):
// \pc_next[20]~84_combout  = (\pc[22]~34_combout  & ((\pc_next[20]~83_combout  & (Result_EX_20)) # (!\pc_next[20]~83_combout  & ((\input_a~158_combout ))))) # (!\pc[22]~34_combout  & (\pc_next[20]~83_combout ))

	.dataa(\pc[22]~34_combout ),
	.datab(\pc_next[20]~83_combout ),
	.datac(Result_EX_20),
	.datad(\input_a~158_combout ),
	.cin(gnd),
	.combout(\pc_next[20]~84_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~84 .lut_mask = 16'hE6C4;
defparam \pc_next[20]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N26
cycloneive_lcell_comb \pc_next[20]~85 (
// Equation(s):
// \pc_next[20]~85_combout  = (\pc[22]~28_combout  & (\pc_next_branch[20]~36_combout )) # (!\pc[22]~28_combout  & ((\pc_next[20]~84_combout )))

	.dataa(\pc_next_branch[20]~36_combout ),
	.datab(\pc[22]~28_combout ),
	.datac(gnd),
	.datad(\pc_next[20]~84_combout ),
	.cin(gnd),
	.combout(\pc_next[20]~85_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~85 .lut_mask = 16'hBB88;
defparam \pc_next[20]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N18
cycloneive_lcell_comb \pc_next[20]~86 (
// Equation(s):
// \pc_next[20]~86_combout  = (\pc_next[20]~85_combout  & (((!\pc[1]~26_combout  & \pc_next_plus4[20]~36_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[20]~85_combout  & (!\pc[1]~26_combout  & ((\pc_next_plus4[20]~36_combout ))))

	.dataa(\pc_next[20]~85_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next[27]~9_combout ),
	.datad(\pc_next_plus4[20]~36_combout ),
	.cin(gnd),
	.combout(\pc_next[20]~86_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~86 .lut_mask = 16'h3B0A;
defparam \pc_next[20]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N2
cycloneive_lcell_comb \input_a~159 (
// Equation(s):
// \input_a~159_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_23)) # (!MemToReg_MEM1 & ((CalcData_MEM_23)))))

	.dataa(\PR|ReadData_MEM [23]),
	.datab(\PR|CalcData_MEM [23]),
	.datac(\PR|MemToReg_MEM~q ),
	.datad(\Equal24~0_combout ),
	.cin(gnd),
	.combout(\input_a~159_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~159 .lut_mask = 16'hAC00;
defparam \input_a~159 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \pc_next[23]~87 (
// Equation(s):
// \pc_next[23]~87_combout  = (\pc[22]~38_combout  & (((\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & ((\input_a~159_combout ))) # (!\pc[22]~34_combout  & (ALUSrc1_ID_23))))

	.dataa(\pc[22]~38_combout ),
	.datab(\PR|ALUSrc1_ID [23]),
	.datac(\pc[22]~34_combout ),
	.datad(\input_a~159_combout ),
	.cin(gnd),
	.combout(\pc_next[23]~87_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~87 .lut_mask = 16'hF4A4;
defparam \pc_next[23]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \pc_next[23]~88 (
// Equation(s):
// \pc_next[23]~88_combout  = (\pc[22]~38_combout  & ((\pc_next[23]~87_combout  & (Result_EX_23)) # (!\pc_next[23]~87_combout  & ((Instr_ID_21))))) # (!\pc[22]~38_combout  & (\pc_next[23]~87_combout ))

	.dataa(\pc[22]~38_combout ),
	.datab(\pc_next[23]~87_combout ),
	.datac(Result_EX_23),
	.datad(\PR|Instr_ID [21]),
	.cin(gnd),
	.combout(\pc_next[23]~88_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~88 .lut_mask = 16'hE6C4;
defparam \pc_next[23]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N10
cycloneive_lcell_comb \pc_next_branch[22]~40 (
// Equation(s):
// \pc_next_branch[22]~40_combout  = ((nextPC_ID_22 $ (Instr_ID_15 $ (!\pc_next_branch[21]~39 )))) # (GND)
// \pc_next_branch[22]~41  = CARRY((nextPC_ID_22 & ((Instr_ID_15) # (!\pc_next_branch[21]~39 ))) # (!nextPC_ID_22 & (Instr_ID_15 & !\pc_next_branch[21]~39 )))

	.dataa(\PR|nextPC_ID [22]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[21]~39 ),
	.combout(\pc_next_branch[22]~40_combout ),
	.cout(\pc_next_branch[22]~41 ));
// synopsys translate_off
defparam \pc_next_branch[22]~40 .lut_mask = 16'h698E;
defparam \pc_next_branch[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \pc_next_branch[23]~42 (
// Equation(s):
// \pc_next_branch[23]~42_combout  = (Instr_ID_15 & ((nextPC_ID_23 & (\pc_next_branch[22]~41  & VCC)) # (!nextPC_ID_23 & (!\pc_next_branch[22]~41 )))) # (!Instr_ID_15 & ((nextPC_ID_23 & (!\pc_next_branch[22]~41 )) # (!nextPC_ID_23 & ((\pc_next_branch[22]~41 
// ) # (GND)))))
// \pc_next_branch[23]~43  = CARRY((Instr_ID_15 & (!nextPC_ID_23 & !\pc_next_branch[22]~41 )) # (!Instr_ID_15 & ((!\pc_next_branch[22]~41 ) # (!nextPC_ID_23))))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [23]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[22]~41 ),
	.combout(\pc_next_branch[23]~42_combout ),
	.cout(\pc_next_branch[23]~43 ));
// synopsys translate_off
defparam \pc_next_branch[23]~42 .lut_mask = 16'h9617;
defparam \pc_next_branch[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N26
cycloneive_lcell_comb \pc_next[23]~89 (
// Equation(s):
// \pc_next[23]~89_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[23]~42_combout ))) # (!\pc[22]~28_combout  & (\pc_next[23]~88_combout ))

	.dataa(gnd),
	.datab(\pc_next[23]~88_combout ),
	.datac(\pc_next_branch[23]~42_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[23]~89_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~89 .lut_mask = 16'hF0CC;
defparam \pc_next[23]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N10
cycloneive_lcell_comb \pc_next_plus4[22]~40 (
// Equation(s):
// \pc_next_plus4[22]~40_combout  = (pc_22 & (\pc_next_plus4[21]~39  $ (GND))) # (!pc_22 & (!\pc_next_plus4[21]~39  & VCC))
// \pc_next_plus4[22]~41  = CARRY((pc_22 & !\pc_next_plus4[21]~39 ))

	.dataa(pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[21]~39 ),
	.combout(\pc_next_plus4[22]~40_combout ),
	.cout(\pc_next_plus4[22]~41 ));
// synopsys translate_off
defparam \pc_next_plus4[22]~40 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N12
cycloneive_lcell_comb \pc_next_plus4[23]~42 (
// Equation(s):
// \pc_next_plus4[23]~42_combout  = (pc_23 & (!\pc_next_plus4[22]~41 )) # (!pc_23 & ((\pc_next_plus4[22]~41 ) # (GND)))
// \pc_next_plus4[23]~43  = CARRY((!\pc_next_plus4[22]~41 ) # (!pc_23))

	.dataa(pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[22]~41 ),
	.combout(\pc_next_plus4[23]~42_combout ),
	.cout(\pc_next_plus4[23]~43 ));
// synopsys translate_off
defparam \pc_next_plus4[23]~42 .lut_mask = 16'h5A5F;
defparam \pc_next_plus4[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N12
cycloneive_lcell_comb \pc_next[23]~90 (
// Equation(s):
// \pc_next[23]~90_combout  = (\pc_next[23]~89_combout  & (((\pc_next_plus4[23]~42_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[23]~89_combout  & (((\pc_next_plus4[23]~42_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[23]~89_combout ),
	.datab(\pc_next[27]~9_combout ),
	.datac(\pc_next_plus4[23]~42_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[23]~90_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~90 .lut_mask = 16'h22F2;
defparam \pc_next[23]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \input_a~160 (
// Equation(s):
// \input_a~160_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_22))) # (!MemToReg_MEM1 & (CalcData_MEM_22))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|CalcData_MEM [22]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|ReadData_MEM [22]),
	.cin(gnd),
	.combout(\input_a~160_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~160 .lut_mask = 16'hE040;
defparam \input_a~160 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \pc_next[22]~91 (
// Equation(s):
// \pc_next[22]~91_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & ((Instr_ID_20))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_22))))

	.dataa(\pc[22]~34_combout ),
	.datab(\PR|ALUSrc1_ID [22]),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [20]),
	.cin(gnd),
	.combout(\pc_next[22]~91_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~91 .lut_mask = 16'hF4A4;
defparam \pc_next[22]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \pc_next[22]~92 (
// Equation(s):
// \pc_next[22]~92_combout  = (\pc[22]~34_combout  & ((\pc_next[22]~91_combout  & ((Result_EX_22))) # (!\pc_next[22]~91_combout  & (\input_a~160_combout )))) # (!\pc[22]~34_combout  & (((\pc_next[22]~91_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(\input_a~160_combout ),
	.datac(\pc_next[22]~91_combout ),
	.datad(Result_EX_22),
	.cin(gnd),
	.combout(\pc_next[22]~92_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~92 .lut_mask = 16'hF858;
defparam \pc_next[22]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N10
cycloneive_lcell_comb \pc_next[22]~93 (
// Equation(s):
// \pc_next[22]~93_combout  = (\pc[22]~28_combout  & (\pc_next_branch[22]~40_combout )) # (!\pc[22]~28_combout  & ((\pc_next[22]~92_combout )))

	.dataa(\pc[22]~28_combout ),
	.datab(\pc_next_branch[22]~40_combout ),
	.datac(gnd),
	.datad(\pc_next[22]~92_combout ),
	.cin(gnd),
	.combout(\pc_next[22]~93_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~93 .lut_mask = 16'hDD88;
defparam \pc_next[22]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N14
cycloneive_lcell_comb \pc_next[22]~94 (
// Equation(s):
// \pc_next[22]~94_combout  = (\pc_next[22]~93_combout  & (((\pc_next_plus4[22]~40_combout  & !\pc[1]~26_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[22]~93_combout  & (((\pc_next_plus4[22]~40_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[22]~93_combout ),
	.datab(\pc_next[27]~9_combout ),
	.datac(\pc_next_plus4[22]~40_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[22]~94_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~94 .lut_mask = 16'h22F2;
defparam \pc_next[22]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N20
cycloneive_lcell_comb \input_a~161 (
// Equation(s):
// \input_a~161_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_25)) # (!MemToReg_MEM1 & ((CalcData_MEM_25)))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [25]),
	.datad(\PR|CalcData_MEM [25]),
	.cin(gnd),
	.combout(\input_a~161_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~161 .lut_mask = 16'hC480;
defparam \input_a~161 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N12
cycloneive_lcell_comb \pc_next[25]~95 (
// Equation(s):
// \pc_next[25]~95_combout  = (\pc[22]~38_combout  & (\pc[22]~34_combout )) # (!\pc[22]~38_combout  & ((\pc[22]~34_combout  & ((\input_a~161_combout ))) # (!\pc[22]~34_combout  & (ALUSrc1_ID_25))))

	.dataa(\pc[22]~38_combout ),
	.datab(\pc[22]~34_combout ),
	.datac(\PR|ALUSrc1_ID [25]),
	.datad(\input_a~161_combout ),
	.cin(gnd),
	.combout(\pc_next[25]~95_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~95 .lut_mask = 16'hDC98;
defparam \pc_next[25]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N28
cycloneive_lcell_comb \pc_next[25]~96 (
// Equation(s):
// \pc_next[25]~96_combout  = (\pc[22]~38_combout  & ((\pc_next[25]~95_combout  & ((Result_EX_25))) # (!\pc_next[25]~95_combout  & (Instr_ID_23)))) # (!\pc[22]~38_combout  & (((\pc_next[25]~95_combout ))))

	.dataa(\pc[22]~38_combout ),
	.datab(\PR|Instr_ID [23]),
	.datac(Result_EX_25),
	.datad(\pc_next[25]~95_combout ),
	.cin(gnd),
	.combout(\pc_next[25]~96_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~96 .lut_mask = 16'hF588;
defparam \pc_next[25]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N14
cycloneive_lcell_comb \pc_next_branch[24]~44 (
// Equation(s):
// \pc_next_branch[24]~44_combout  = ((nextPC_ID_24 $ (Instr_ID_15 $ (!\pc_next_branch[23]~43 )))) # (GND)
// \pc_next_branch[24]~45  = CARRY((nextPC_ID_24 & ((Instr_ID_15) # (!\pc_next_branch[23]~43 ))) # (!nextPC_ID_24 & (Instr_ID_15 & !\pc_next_branch[23]~43 )))

	.dataa(\PR|nextPC_ID [24]),
	.datab(\PR|Instr_ID [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[23]~43 ),
	.combout(\pc_next_branch[24]~44_combout ),
	.cout(\pc_next_branch[24]~45 ));
// synopsys translate_off
defparam \pc_next_branch[24]~44 .lut_mask = 16'h698E;
defparam \pc_next_branch[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N16
cycloneive_lcell_comb \pc_next_branch[25]~46 (
// Equation(s):
// \pc_next_branch[25]~46_combout  = (Instr_ID_15 & ((nextPC_ID_25 & (\pc_next_branch[24]~45  & VCC)) # (!nextPC_ID_25 & (!\pc_next_branch[24]~45 )))) # (!Instr_ID_15 & ((nextPC_ID_25 & (!\pc_next_branch[24]~45 )) # (!nextPC_ID_25 & ((\pc_next_branch[24]~45 
// ) # (GND)))))
// \pc_next_branch[25]~47  = CARRY((Instr_ID_15 & (!nextPC_ID_25 & !\pc_next_branch[24]~45 )) # (!Instr_ID_15 & ((!\pc_next_branch[24]~45 ) # (!nextPC_ID_25))))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [25]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[24]~45 ),
	.combout(\pc_next_branch[25]~46_combout ),
	.cout(\pc_next_branch[25]~47 ));
// synopsys translate_off
defparam \pc_next_branch[25]~46 .lut_mask = 16'h9617;
defparam \pc_next_branch[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \pc_next[25]~97 (
// Equation(s):
// \pc_next[25]~97_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[25]~46_combout ))) # (!\pc[22]~28_combout  & (\pc_next[25]~96_combout ))

	.dataa(\pc[22]~28_combout ),
	.datab(gnd),
	.datac(\pc_next[25]~96_combout ),
	.datad(\pc_next_branch[25]~46_combout ),
	.cin(gnd),
	.combout(\pc_next[25]~97_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~97 .lut_mask = 16'hFA50;
defparam \pc_next[25]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N14
cycloneive_lcell_comb \pc_next_plus4[24]~44 (
// Equation(s):
// \pc_next_plus4[24]~44_combout  = (pc_24 & (\pc_next_plus4[23]~43  $ (GND))) # (!pc_24 & (!\pc_next_plus4[23]~43  & VCC))
// \pc_next_plus4[24]~45  = CARRY((pc_24 & !\pc_next_plus4[23]~43 ))

	.dataa(pc_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[23]~43 ),
	.combout(\pc_next_plus4[24]~44_combout ),
	.cout(\pc_next_plus4[24]~45 ));
// synopsys translate_off
defparam \pc_next_plus4[24]~44 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N16
cycloneive_lcell_comb \pc_next_plus4[25]~46 (
// Equation(s):
// \pc_next_plus4[25]~46_combout  = (pc_25 & (!\pc_next_plus4[24]~45 )) # (!pc_25 & ((\pc_next_plus4[24]~45 ) # (GND)))
// \pc_next_plus4[25]~47  = CARRY((!\pc_next_plus4[24]~45 ) # (!pc_25))

	.dataa(pc_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[24]~45 ),
	.combout(\pc_next_plus4[25]~46_combout ),
	.cout(\pc_next_plus4[25]~47 ));
// synopsys translate_off
defparam \pc_next_plus4[25]~46 .lut_mask = 16'h5A5F;
defparam \pc_next_plus4[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \pc_next[25]~98 (
// Equation(s):
// \pc_next[25]~98_combout  = (\pc_next[25]~97_combout  & (((!\pc[1]~26_combout  & \pc_next_plus4[25]~46_combout )) # (!\pc_next[27]~9_combout ))) # (!\pc_next[25]~97_combout  & (!\pc[1]~26_combout  & (\pc_next_plus4[25]~46_combout )))

	.dataa(\pc_next[25]~97_combout ),
	.datab(\pc[1]~26_combout ),
	.datac(\pc_next_plus4[25]~46_combout ),
	.datad(\pc_next[27]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[25]~98_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~98 .lut_mask = 16'h30BA;
defparam \pc_next[25]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \pc_next[24]~99 (
// Equation(s):
// \pc_next[24]~99_combout  = (\pc[22]~34_combout  & (((\pc[22]~38_combout )))) # (!\pc[22]~34_combout  & ((\pc[22]~38_combout  & ((Instr_ID_22))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_24))))

	.dataa(\PR|ALUSrc1_ID [24]),
	.datab(\pc[22]~34_combout ),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [22]),
	.cin(gnd),
	.combout(\pc_next[24]~99_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~99 .lut_mask = 16'hF2C2;
defparam \pc_next[24]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \pc_next[24]~100 (
// Equation(s):
// \pc_next[24]~100_combout  = (\pc[22]~34_combout  & ((\pc_next[24]~99_combout  & ((Result_EX_24))) # (!\pc_next[24]~99_combout  & (\input_a~162_combout )))) # (!\pc[22]~34_combout  & (((\pc_next[24]~99_combout ))))

	.dataa(\input_a~162_combout ),
	.datab(\pc[22]~34_combout ),
	.datac(Result_EX_24),
	.datad(\pc_next[24]~99_combout ),
	.cin(gnd),
	.combout(\pc_next[24]~100_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~100 .lut_mask = 16'hF388;
defparam \pc_next[24]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \pc_next[24]~101 (
// Equation(s):
// \pc_next[24]~101_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[24]~44_combout ))) # (!\pc[22]~28_combout  & (\pc_next[24]~100_combout ))

	.dataa(gnd),
	.datab(\pc_next[24]~100_combout ),
	.datac(\pc_next_branch[24]~44_combout ),
	.datad(\pc[22]~28_combout ),
	.cin(gnd),
	.combout(\pc_next[24]~101_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~101 .lut_mask = 16'hF0CC;
defparam \pc_next[24]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \pc_next[24]~102 (
// Equation(s):
// \pc_next[24]~102_combout  = (\pc_next[27]~9_combout  & (((\pc_next_plus4[24]~44_combout  & !\pc[1]~26_combout )))) # (!\pc_next[27]~9_combout  & ((\pc_next[24]~101_combout ) # ((\pc_next_plus4[24]~44_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[27]~9_combout ),
	.datab(\pc_next[24]~101_combout ),
	.datac(\pc_next_plus4[24]~44_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[24]~102_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~102 .lut_mask = 16'h44F4;
defparam \pc_next[24]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N18
cycloneive_lcell_comb \pc_next_plus4[26]~48 (
// Equation(s):
// \pc_next_plus4[26]~48_combout  = (pc_26 & (\pc_next_plus4[25]~47  $ (GND))) # (!pc_26 & (!\pc_next_plus4[25]~47  & VCC))
// \pc_next_plus4[26]~49  = CARRY((pc_26 & !\pc_next_plus4[25]~47 ))

	.dataa(pc_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[25]~47 ),
	.combout(\pc_next_plus4[26]~48_combout ),
	.cout(\pc_next_plus4[26]~49 ));
// synopsys translate_off
defparam \pc_next_plus4[26]~48 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N20
cycloneive_lcell_comb \pc_next_plus4[27]~50 (
// Equation(s):
// \pc_next_plus4[27]~50_combout  = (pc_27 & (!\pc_next_plus4[26]~49 )) # (!pc_27 & ((\pc_next_plus4[26]~49 ) # (GND)))
// \pc_next_plus4[27]~51  = CARRY((!\pc_next_plus4[26]~49 ) # (!pc_27))

	.dataa(gnd),
	.datab(pc_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[26]~49 ),
	.combout(\pc_next_plus4[27]~50_combout ),
	.cout(\pc_next_plus4[27]~51 ));
// synopsys translate_off
defparam \pc_next_plus4[27]~50 .lut_mask = 16'h3C3F;
defparam \pc_next_plus4[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \pc_next[27]~104 (
// Equation(s):
// \pc_next[27]~104_combout  = (\pc_next[27]~103_combout  & ((Result_EX_27) # ((!\pc[22]~38_combout )))) # (!\pc_next[27]~103_combout  & (((\pc[22]~38_combout  & Instr_ID_25))))

	.dataa(\pc_next[27]~103_combout ),
	.datab(Result_EX_27),
	.datac(\pc[22]~38_combout ),
	.datad(\PR|Instr_ID [25]),
	.cin(gnd),
	.combout(\pc_next[27]~104_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~104 .lut_mask = 16'hDA8A;
defparam \pc_next[27]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N18
cycloneive_lcell_comb \pc_next_branch[26]~48 (
// Equation(s):
// \pc_next_branch[26]~48_combout  = ((Instr_ID_15 $ (nextPC_ID_26 $ (!\pc_next_branch[25]~47 )))) # (GND)
// \pc_next_branch[26]~49  = CARRY((Instr_ID_15 & ((nextPC_ID_26) # (!\pc_next_branch[25]~47 ))) # (!Instr_ID_15 & (nextPC_ID_26 & !\pc_next_branch[25]~47 )))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [26]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[25]~47 ),
	.combout(\pc_next_branch[26]~48_combout ),
	.cout(\pc_next_branch[26]~49 ));
// synopsys translate_off
defparam \pc_next_branch[26]~48 .lut_mask = 16'h698E;
defparam \pc_next_branch[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N20
cycloneive_lcell_comb \pc_next_branch[27]~50 (
// Equation(s):
// \pc_next_branch[27]~50_combout  = (Instr_ID_15 & ((nextPC_ID_27 & (\pc_next_branch[26]~49  & VCC)) # (!nextPC_ID_27 & (!\pc_next_branch[26]~49 )))) # (!Instr_ID_15 & ((nextPC_ID_27 & (!\pc_next_branch[26]~49 )) # (!nextPC_ID_27 & ((\pc_next_branch[26]~49 
// ) # (GND)))))
// \pc_next_branch[27]~51  = CARRY((Instr_ID_15 & (!nextPC_ID_27 & !\pc_next_branch[26]~49 )) # (!Instr_ID_15 & ((!\pc_next_branch[26]~49 ) # (!nextPC_ID_27))))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [27]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[26]~49 ),
	.combout(\pc_next_branch[27]~50_combout ),
	.cout(\pc_next_branch[27]~51 ));
// synopsys translate_off
defparam \pc_next_branch[27]~50 .lut_mask = 16'h9617;
defparam \pc_next_branch[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \pc_next[27]~105 (
// Equation(s):
// \pc_next[27]~105_combout  = (\pc[22]~28_combout  & ((\pc_next_branch[27]~50_combout ))) # (!\pc[22]~28_combout  & (\pc_next[27]~104_combout ))

	.dataa(\pc[22]~28_combout ),
	.datab(\pc_next[27]~104_combout ),
	.datac(\pc_next_branch[27]~50_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_next[27]~105_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~105 .lut_mask = 16'hE4E4;
defparam \pc_next[27]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \pc_next[27]~106 (
// Equation(s):
// \pc_next[27]~106_combout  = (\pc_next[27]~9_combout  & (\pc_next_plus4[27]~50_combout  & ((!\pc[1]~26_combout )))) # (!\pc_next[27]~9_combout  & ((\pc_next[27]~105_combout ) # ((\pc_next_plus4[27]~50_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[27]~9_combout ),
	.datab(\pc_next_plus4[27]~50_combout ),
	.datac(\pc_next[27]~105_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[27]~106_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~106 .lut_mask = 16'h50DC;
defparam \pc_next[27]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \input_a~164 (
// Equation(s):
// \input_a~164_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_26))) # (!MemToReg_MEM1 & (CalcData_MEM_26))))

	.dataa(\PR|CalcData_MEM [26]),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [26]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~164_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~164 .lut_mask = 16'hC088;
defparam \input_a~164 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \pc_next[26]~107 (
// Equation(s):
// \pc_next[26]~107_combout  = (\pc[22]~38_combout  & (((Instr_ID_24) # (\pc[22]~34_combout )))) # (!\pc[22]~38_combout  & (ALUSrc1_ID_26 & ((!\pc[22]~34_combout ))))

	.dataa(\PR|ALUSrc1_ID [26]),
	.datab(\PR|Instr_ID [24]),
	.datac(\pc[22]~38_combout ),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~107_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~107 .lut_mask = 16'hF0CA;
defparam \pc_next[26]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \pc_next[26]~108 (
// Equation(s):
// \pc_next[26]~108_combout  = (\pc[22]~34_combout  & ((\pc_next[26]~107_combout  & (Result_EX_26)) # (!\pc_next[26]~107_combout  & ((\input_a~164_combout ))))) # (!\pc[22]~34_combout  & (((\pc_next[26]~107_combout ))))

	.dataa(\pc[22]~34_combout ),
	.datab(Result_EX_26),
	.datac(\input_a~164_combout ),
	.datad(\pc_next[26]~107_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~108_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~108 .lut_mask = 16'hDDA0;
defparam \pc_next[26]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N24
cycloneive_lcell_comb \pc_next[26]~109 (
// Equation(s):
// \pc_next[26]~109_combout  = (\pc[22]~28_combout  & (\pc_next_branch[26]~48_combout )) # (!\pc[22]~28_combout  & ((\pc_next[26]~108_combout )))

	.dataa(\pc[22]~28_combout ),
	.datab(\pc_next_branch[26]~48_combout ),
	.datac(\pc_next[26]~108_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_next[26]~109_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~109 .lut_mask = 16'hD8D8;
defparam \pc_next[26]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \pc_next[26]~110 (
// Equation(s):
// \pc_next[26]~110_combout  = (\pc_next[27]~9_combout  & (\pc_next_plus4[26]~48_combout  & ((!\pc[1]~26_combout )))) # (!\pc_next[27]~9_combout  & ((\pc_next[26]~109_combout ) # ((\pc_next_plus4[26]~48_combout  & !\pc[1]~26_combout ))))

	.dataa(\pc_next[27]~9_combout ),
	.datab(\pc_next_plus4[26]~48_combout ),
	.datac(\pc_next[26]~109_combout ),
	.datad(\pc[1]~26_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~110_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~110 .lut_mask = 16'h50DC;
defparam \pc_next[26]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \pc[29]~35 (
// Equation(s):
// \pc[29]~35_combout  = (jump_ID_2) # ((jump_ID_0) # ((!always03 & !src1_hazard_t)))

	.dataa(\HZ|always0~8_combout ),
	.datab(\PR|jump_ID [2]),
	.datac(\PR|jump_ID [0]),
	.datad(\HZ|src1_hazard_t~1_combout ),
	.cin(gnd),
	.combout(\pc[29]~35_combout ),
	.cout());
// synopsys translate_off
defparam \pc[29]~35 .lut_mask = 16'hFCFD;
defparam \pc[29]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N18
cycloneive_lcell_comb \Equal23~0 (
// Equation(s):
// \Equal23~0_combout  = (!MemToReg_EX1 & always03)

	.dataa(gnd),
	.datab(MemToReg_EX),
	.datac(\HZ|always0~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal23~0 .lut_mask = 16'h3030;
defparam \Equal23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N30
cycloneive_lcell_comb \pc[29]~31 (
// Equation(s):
// \pc[29]~31_combout  = (jump_ID_2 & ((\pc[29]~35_combout  & (!\pc[29]~29_combout )) # (!\pc[29]~35_combout  & ((!\Equal23~0_combout )))))

	.dataa(\pc[29]~29_combout ),
	.datab(\pc[29]~35_combout ),
	.datac(\PR|jump_ID [2]),
	.datad(\Equal23~0_combout ),
	.cin(gnd),
	.combout(\pc[29]~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc[29]~31 .lut_mask = 16'h4070;
defparam \pc[29]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N20
cycloneive_lcell_comb \pc[29]~30 (
// Equation(s):
// \pc[29]~30_combout  = (jump_ID_2 & (\pc[29]~29_combout )) # (!jump_ID_2 & ((\pc[22]~34_combout  & ((\Equal23~0_combout ))) # (!\pc[22]~34_combout  & (\pc[29]~29_combout ))))

	.dataa(\pc[29]~29_combout ),
	.datab(\Equal23~0_combout ),
	.datac(\PR|jump_ID [2]),
	.datad(\pc[22]~34_combout ),
	.cin(gnd),
	.combout(\pc[29]~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc[29]~30 .lut_mask = 16'hACAA;
defparam \pc[29]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N8
cycloneive_lcell_comb \pc_next[29]~111 (
// Equation(s):
// \pc_next[29]~111_combout  = (\pc[29]~30_combout  & (((Result_EX_29) # (\pc[29]~35_combout )))) # (!\pc[29]~30_combout  & (\input_a~165_combout  & ((!\pc[29]~35_combout ))))

	.dataa(\input_a~165_combout ),
	.datab(Result_EX_29),
	.datac(\pc[29]~30_combout ),
	.datad(\pc[29]~35_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~111_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~111 .lut_mask = 16'hF0CA;
defparam \pc_next[29]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N22
cycloneive_lcell_comb \pc_next_branch[28]~52 (
// Equation(s):
// \pc_next_branch[28]~52_combout  = ((Instr_ID_15 $ (nextPC_ID_28 $ (!\pc_next_branch[27]~51 )))) # (GND)
// \pc_next_branch[28]~53  = CARRY((Instr_ID_15 & ((nextPC_ID_28) # (!\pc_next_branch[27]~51 ))) # (!Instr_ID_15 & (nextPC_ID_28 & !\pc_next_branch[27]~51 )))

	.dataa(\PR|Instr_ID [15]),
	.datab(\PR|nextPC_ID [28]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_branch[27]~51 ),
	.combout(\pc_next_branch[28]~52_combout ),
	.cout(\pc_next_branch[28]~53 ));
// synopsys translate_off
defparam \pc_next_branch[28]~52 .lut_mask = 16'h698E;
defparam \pc_next_branch[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N14
cycloneive_lcell_comb \pc_next[29]~112 (
// Equation(s):
// \pc_next[29]~112_combout  = (\pc[29]~35_combout  & ((\pc_next[29]~111_combout  & ((\pc_next_branch[29]~54_combout ))) # (!\pc_next[29]~111_combout  & (ALUSrc1_ID_29)))) # (!\pc[29]~35_combout  & (((\pc_next[29]~111_combout ))))

	.dataa(\pc[29]~35_combout ),
	.datab(\PR|ALUSrc1_ID [29]),
	.datac(\pc_next[29]~111_combout ),
	.datad(\pc_next_branch[29]~54_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~112_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~112 .lut_mask = 16'hF858;
defparam \pc_next[29]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N22
cycloneive_lcell_comb \pc_next_plus4[28]~52 (
// Equation(s):
// \pc_next_plus4[28]~52_combout  = (pc_28 & (\pc_next_plus4[27]~51  $ (GND))) # (!pc_28 & (!\pc_next_plus4[27]~51  & VCC))
// \pc_next_plus4[28]~53  = CARRY((pc_28 & !\pc_next_plus4[27]~51 ))

	.dataa(pc_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[27]~51 ),
	.combout(\pc_next_plus4[28]~52_combout ),
	.cout(\pc_next_plus4[28]~53 ));
// synopsys translate_off
defparam \pc_next_plus4[28]~52 .lut_mask = 16'hA50A;
defparam \pc_next_plus4[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N24
cycloneive_lcell_comb \pc_next_plus4[29]~54 (
// Equation(s):
// \pc_next_plus4[29]~54_combout  = (pc_29 & (!\pc_next_plus4[28]~53 )) # (!pc_29 & ((\pc_next_plus4[28]~53 ) # (GND)))
// \pc_next_plus4[29]~55  = CARRY((!\pc_next_plus4[28]~53 ) # (!pc_29))

	.dataa(pc_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[28]~53 ),
	.combout(\pc_next_plus4[29]~54_combout ),
	.cout(\pc_next_plus4[29]~55 ));
// synopsys translate_off
defparam \pc_next_plus4[29]~54 .lut_mask = 16'h5A5F;
defparam \pc_next_plus4[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \pc[29]~36 (
// Equation(s):
// \pc[29]~36_combout  = (jump_ID_0 & (((jump_ID_2) # (Equal11)))) # (!jump_ID_0 & ((jump_ID_1) # ((jump_ID_2 & !Equal11))))

	.dataa(\PR|jump_ID [1]),
	.datab(\PR|jump_ID [2]),
	.datac(\PR|jump_ID [0]),
	.datad(\ALU|Equal11~11_combout ),
	.cin(gnd),
	.combout(\pc[29]~36_combout ),
	.cout());
// synopsys translate_off
defparam \pc[29]~36 .lut_mask = 16'hFACE;
defparam \pc[29]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \pc_next[29]~113 (
// Equation(s):
// \pc_next[29]~113_combout  = (\pc[29]~36_combout  & (!\pc[29]~31_combout  & (\pc_next[29]~112_combout ))) # (!\pc[29]~36_combout  & (((\pc_next_plus4[29]~54_combout ))))

	.dataa(\pc[29]~31_combout ),
	.datab(\pc_next[29]~112_combout ),
	.datac(\pc_next_plus4[29]~54_combout ),
	.datad(\pc[29]~36_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~113_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~113 .lut_mask = 16'h44F0;
defparam \pc_next[29]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \pc[31]~32 (
// Equation(s):
// \pc[31]~32_combout  = (!\Equal8~0_combout  & (always1 & ((\branch~0_combout ) # (!always0))))

	.dataa(\Equal8~0_combout ),
	.datab(always1),
	.datac(always0),
	.datad(\branch~0_combout ),
	.cin(gnd),
	.combout(\pc[31]~32_combout ),
	.cout());
// synopsys translate_off
defparam \pc[31]~32 .lut_mask = 16'h4404;
defparam \pc[31]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N18
cycloneive_lcell_comb \pc_next[28]~115 (
// Equation(s):
// \pc_next[28]~115_combout  = (\pc_next[28]~114_combout  & (((\pc_next_branch[28]~52_combout ) # (!\pc[29]~30_combout )))) # (!\pc_next[28]~114_combout  & (Result_EX_28 & (\pc[29]~30_combout )))

	.dataa(\pc_next[28]~114_combout ),
	.datab(Result_EX_28),
	.datac(\pc[29]~30_combout ),
	.datad(\pc_next_branch[28]~52_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~115_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~115 .lut_mask = 16'hEA4A;
defparam \pc_next[28]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N2
cycloneive_lcell_comb \pc_next[28]~116 (
// Equation(s):
// \pc_next[28]~116_combout  = (\pc[29]~36_combout  & (!\pc[29]~31_combout  & ((\pc_next[28]~115_combout )))) # (!\pc[29]~36_combout  & (((\pc_next_plus4[28]~52_combout ))))

	.dataa(\pc[29]~31_combout ),
	.datab(\pc_next_plus4[28]~52_combout ),
	.datac(\pc_next[28]~115_combout ),
	.datad(\pc[29]~36_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~116_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~116 .lut_mask = 16'h50CC;
defparam \pc_next[28]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \input_a~167 (
// Equation(s):
// \input_a~167_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & ((ReadData_MEM_31))) # (!MemToReg_MEM1 & (CalcData_MEM_31))))

	.dataa(\PR|CalcData_MEM [31]),
	.datab(\Equal24~0_combout ),
	.datac(\PR|ReadData_MEM [31]),
	.datad(\PR|MemToReg_MEM~q ),
	.cin(gnd),
	.combout(\input_a~167_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~167 .lut_mask = 16'hC088;
defparam \input_a~167 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N4
cycloneive_lcell_comb \pc_next[31]~117 (
// Equation(s):
// \pc_next[31]~117_combout  = (\pc[29]~30_combout  & ((Result_EX_31) # ((\pc[29]~35_combout )))) # (!\pc[29]~30_combout  & (((\input_a~167_combout  & !\pc[29]~35_combout ))))

	.dataa(\pc[29]~30_combout ),
	.datab(Result_EX_31),
	.datac(\input_a~167_combout ),
	.datad(\pc[29]~35_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~117_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~117 .lut_mask = 16'hAAD8;
defparam \pc_next[31]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N2
cycloneive_lcell_comb \pc_next[31]~118 (
// Equation(s):
// \pc_next[31]~118_combout  = (\pc_next[31]~117_combout  & ((\pc_next_branch[31]~58_combout ) # ((!\pc[29]~35_combout )))) # (!\pc_next[31]~117_combout  & (((ALUSrc1_ID_31 & \pc[29]~35_combout ))))

	.dataa(\pc_next_branch[31]~58_combout ),
	.datab(\PR|ALUSrc1_ID [31]),
	.datac(\pc_next[31]~117_combout ),
	.datad(\pc[29]~35_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~118_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~118 .lut_mask = 16'hACF0;
defparam \pc_next[31]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N26
cycloneive_lcell_comb \pc_next_plus4[30]~56 (
// Equation(s):
// \pc_next_plus4[30]~56_combout  = (pc_30 & (\pc_next_plus4[29]~55  $ (GND))) # (!pc_30 & (!\pc_next_plus4[29]~55  & VCC))
// \pc_next_plus4[30]~57  = CARRY((pc_30 & !\pc_next_plus4[29]~55 ))

	.dataa(gnd),
	.datab(pc_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_next_plus4[29]~55 ),
	.combout(\pc_next_plus4[30]~56_combout ),
	.cout(\pc_next_plus4[30]~57 ));
// synopsys translate_off
defparam \pc_next_plus4[30]~56 .lut_mask = 16'hC30C;
defparam \pc_next_plus4[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N28
cycloneive_lcell_comb \pc_next_plus4[31]~58 (
// Equation(s):
// \pc_next_plus4[31]~58_combout  = \pc_next_plus4[30]~57  $ (pc_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_31),
	.cin(\pc_next_plus4[30]~57 ),
	.combout(\pc_next_plus4[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next_plus4[31]~58 .lut_mask = 16'h0FF0;
defparam \pc_next_plus4[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \pc_next[31]~119 (
// Equation(s):
// \pc_next[31]~119_combout  = (\pc[29]~36_combout  & (!\pc[29]~31_combout  & (\pc_next[31]~118_combout ))) # (!\pc[29]~36_combout  & (((\pc_next_plus4[31]~58_combout ))))

	.dataa(\pc[29]~31_combout ),
	.datab(\pc_next[31]~118_combout ),
	.datac(\pc_next_plus4[31]~58_combout ),
	.datad(\pc[29]~36_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~119_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~119 .lut_mask = 16'h44F0;
defparam \pc_next[31]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \input_a~168 (
// Equation(s):
// \input_a~168_combout  = (\Equal24~0_combout  & ((MemToReg_MEM1 & (ReadData_MEM_30)) # (!MemToReg_MEM1 & ((CalcData_MEM_30)))))

	.dataa(\PR|MemToReg_MEM~q ),
	.datab(\PR|ReadData_MEM [30]),
	.datac(\Equal24~0_combout ),
	.datad(\PR|CalcData_MEM [30]),
	.cin(gnd),
	.combout(\input_a~168_combout ),
	.cout());
// synopsys translate_off
defparam \input_a~168 .lut_mask = 16'hD080;
defparam \input_a~168 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N20
cycloneive_lcell_comb \pc_next[30]~120 (
// Equation(s):
// \pc_next[30]~120_combout  = (\pc[29]~30_combout  & (((\pc[29]~35_combout )))) # (!\pc[29]~30_combout  & ((\pc[29]~35_combout  & ((ALUSrc1_ID_30))) # (!\pc[29]~35_combout  & (\input_a~168_combout ))))

	.dataa(\pc[29]~30_combout ),
	.datab(\input_a~168_combout ),
	.datac(\PR|ALUSrc1_ID [30]),
	.datad(\pc[29]~35_combout ),
	.cin(gnd),
	.combout(\pc_next[30]~120_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~120 .lut_mask = 16'hFA44;
defparam \pc_next[30]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N26
cycloneive_lcell_comb \pc_next[30]~121 (
// Equation(s):
// \pc_next[30]~121_combout  = (\pc[29]~30_combout  & ((\pc_next[30]~120_combout  & (\pc_next_branch[30]~56_combout )) # (!\pc_next[30]~120_combout  & ((Result_EX_30))))) # (!\pc[29]~30_combout  & (((\pc_next[30]~120_combout ))))

	.dataa(\pc_next_branch[30]~56_combout ),
	.datab(Result_EX_30),
	.datac(\pc[29]~30_combout ),
	.datad(\pc_next[30]~120_combout ),
	.cin(gnd),
	.combout(\pc_next[30]~121_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~121 .lut_mask = 16'hAFC0;
defparam \pc_next[30]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \pc_next[30]~122 (
// Equation(s):
// \pc_next[30]~122_combout  = (\pc[29]~36_combout  & (\pc_next[30]~121_combout  & ((!\pc[29]~31_combout )))) # (!\pc[29]~36_combout  & (((\pc_next_plus4[30]~56_combout ))))

	.dataa(\pc[29]~36_combout ),
	.datab(\pc_next[30]~121_combout ),
	.datac(\pc_next_plus4[30]~56_combout ),
	.datad(\pc[29]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[30]~122_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~122 .lut_mask = 16'h50D8;
defparam \pc_next[30]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N17
dffeas \halt_reg~_Duplicate_1 (
	.clk(!CLK),
	.d(\halt_reg~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\halt_reg~_Duplicate_1_q ),
	.prn(vcc));
// synopsys translate_off
defparam \halt_reg~_Duplicate_1 .is_wysiwyg = "true";
defparam \halt_reg~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N22
cycloneive_lcell_comb \halt_reg~0 (
// Equation(s):
// \halt_reg~0_combout  = (\halt_reg~_Duplicate_1_q ) # ((halt_MEM1 & !care_ID1))

	.dataa(gnd),
	.datab(\halt_reg~_Duplicate_1_q ),
	.datac(\PR|halt_MEM~q ),
	.datad(\PR|care_ID~q ),
	.cin(gnd),
	.combout(\halt_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~0 .lut_mask = 16'hCCFC;
defparam \halt_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N12
cycloneive_lcell_comb \halt_reg~1 (
// Equation(s):
// \halt_reg~1_combout  = (!ALUOP_ID_2 & (care_ID1 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(\PR|ALUOP_ID [2]),
	.datab(\PR|care_ID~q ),
	.datac(\PR|ALUOP_ID [1]),
	.datad(\PR|ALUOP_ID [3]),
	.cin(gnd),
	.combout(\halt_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~1 .lut_mask = 16'h0040;
defparam \halt_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N30
cycloneive_lcell_comb \halt_reg~2 (
// Equation(s):
// \halt_reg~2_combout  = (ALUOP_ID_0 & (out & (\input_a~61_combout  $ (Add1))))

	.dataa(\input_a~61_combout ),
	.datab(\PR|ALUOP_ID [0]),
	.datac(\ALU|out~0_combout ),
	.datad(\ALU|Add1~62_combout ),
	.cin(gnd),
	.combout(\halt_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~2 .lut_mask = 16'h4080;
defparam \halt_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N8
cycloneive_lcell_comb \halt_reg~3 (
// Equation(s):
// \halt_reg~3_combout  = (!out & !ALUOP_ID_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|out~0_combout ),
	.datad(\PR|ALUOP_ID [0]),
	.cin(gnd),
	.combout(\halt_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~3 .lut_mask = 16'h000F;
defparam \halt_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N0
cycloneive_lcell_comb \halt_reg~4 (
// Equation(s):
// \halt_reg~4_combout  = (Add0) # ((Add03) # ((Add01) # (Add04)))

	.dataa(\ALU|Add0~42_combout ),
	.datab(\ALU|Add0~48_combout ),
	.datac(\ALU|Add0~44_combout ),
	.datad(\ALU|Add0~50_combout ),
	.cin(gnd),
	.combout(\halt_reg~4_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~4 .lut_mask = 16'hFFFE;
defparam \halt_reg~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N26
cycloneive_lcell_comb \halt_reg~5 (
// Equation(s):
// \halt_reg~5_combout  = (Add07) # ((Add09) # (\halt_reg~4_combout ))

	.dataa(gnd),
	.datab(\ALU|Add0~56_combout ),
	.datac(\ALU|Add0~60_combout ),
	.datad(\halt_reg~4_combout ),
	.cin(gnd),
	.combout(\halt_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~5 .lut_mask = 16'hFFFC;
defparam \halt_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N24
cycloneive_lcell_comb \halt_reg~6 (
// Equation(s):
// \halt_reg~6_combout  = (Add02) # ((Equal0) # ((!Equal02) # (!Equal01)))

	.dataa(\ALU|Add0~46_combout ),
	.datab(\ALU|Equal0~0_combout ),
	.datac(\ALU|Equal0~5_combout ),
	.datad(\ALU|Equal0~6_combout ),
	.cin(gnd),
	.combout(\halt_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~6 .lut_mask = 16'hEFFF;
defparam \halt_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N6
cycloneive_lcell_comb \halt_reg~7 (
// Equation(s):
// \halt_reg~7_combout  = (Add05) # ((Add06) # ((Add08) # (\halt_reg~6_combout )))

	.dataa(\ALU|Add0~52_combout ),
	.datab(\ALU|Add0~54_combout ),
	.datac(\ALU|Add0~58_combout ),
	.datad(\halt_reg~6_combout ),
	.cin(gnd),
	.combout(\halt_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~7 .lut_mask = 16'hFFFE;
defparam \halt_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N20
cycloneive_lcell_comb \halt_reg~8 (
// Equation(s):
// \halt_reg~8_combout  = (\halt_reg~3_combout  & ((Add010) # ((\halt_reg~5_combout ) # (\halt_reg~7_combout ))))

	.dataa(\ALU|Add0~62_combout ),
	.datab(\halt_reg~3_combout ),
	.datac(\halt_reg~5_combout ),
	.datad(\halt_reg~7_combout ),
	.cin(gnd),
	.combout(\halt_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~8 .lut_mask = 16'hCCC8;
defparam \halt_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N16
cycloneive_lcell_comb \halt_reg~9 (
// Equation(s):
// \halt_reg~9_combout  = (\halt_reg~0_combout ) # ((\halt_reg~1_combout  & ((\halt_reg~2_combout ) # (\halt_reg~8_combout ))))

	.dataa(\halt_reg~0_combout ),
	.datab(\halt_reg~1_combout ),
	.datac(\halt_reg~2_combout ),
	.datad(\halt_reg~8_combout ),
	.cin(gnd),
	.combout(\halt_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \halt_reg~9 .lut_mask = 16'hEEEA;
defparam \halt_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu_file (
	Add1,
	Add0,
	Add01,
	Add02,
	Add03,
	Add04,
	Add05,
	Add06,
	Add07,
	Add08,
	Add09,
	Add010,
	Result_EX_1,
	Result_EX_0,
	Result_EX_3,
	Result_EX_2,
	Result_EX_4,
	Result_EX_7,
	Result_EX_31,
	ALUOP_ID_1,
	ALUOP_ID_3,
	ALUOP_ID_2,
	input_b,
	input_b1,
	input_a,
	out,
	ALUOP_ID_0,
	input_b2,
	input_a1,
	input_b3,
	input_a2,
	input_b4,
	input_a3,
	input_b5,
	input_a4,
	input_b6,
	input_a5,
	input_b7,
	input_a6,
	input_b8,
	input_a7,
	input_b9,
	input_a8,
	input_b10,
	input_a9,
	input_b11,
	input_a10,
	input_b12,
	input_a11,
	input_b13,
	input_a12,
	input_b14,
	input_a13,
	input_b15,
	input_a14,
	input_b16,
	input_a15,
	input_b17,
	input_a16,
	input_b18,
	input_a17,
	input_b19,
	input_b20,
	input_a18,
	input_b21,
	input_a19,
	input_b22,
	input_a20,
	input_b23,
	input_a21,
	input_b24,
	input_a22,
	input_b25,
	input_a23,
	input_b26,
	input_b27,
	input_a24,
	input_b28,
	input_a25,
	input_b29,
	input_a26,
	input_b30,
	input_b31,
	input_a27,
	input_b32,
	input_b33,
	input_a28,
	input_b34,
	input_b35,
	input_a29,
	input_b36,
	input_b37,
	input_a30,
	input_b38,
	input_b39,
	input_a31,
	Equal0,
	Equal01,
	Equal02,
	Selector30,
	halt_reg,
	Selector28,
	Selector3,
	Selector22,
	Selector2,
	Selector27,
	Selector25,
	input_b40,
	Selector24,
	Selector26,
	Selector4,
	Selector16,
	Selector7,
	Selector6,
	Selector29,
	Selector15,
	Selector5,
	Selector31,
	Selector11,
	Selector10,
	Selector21,
	Selector20,
	Selector9,
	Selector8,
	Selector14,
	Selector13,
	Selector12,
	Selector23,
	Selector19,
	Selector18,
	Selector17,
	Selector0,
	Selector1,
	Equal11,
	devpor,
	devclrn,
	devoe);
output 	Add1;
output 	Add0;
output 	Add01;
output 	Add02;
output 	Add03;
output 	Add04;
output 	Add05;
output 	Add06;
output 	Add07;
output 	Add08;
output 	Add09;
output 	Add010;
input 	Result_EX_1;
input 	Result_EX_0;
input 	Result_EX_3;
input 	Result_EX_2;
input 	Result_EX_4;
input 	Result_EX_7;
input 	Result_EX_31;
input 	ALUOP_ID_1;
input 	ALUOP_ID_3;
input 	ALUOP_ID_2;
input 	input_b;
input 	input_b1;
input 	input_a;
output 	out;
input 	ALUOP_ID_0;
input 	input_b2;
input 	input_a1;
input 	input_b3;
input 	input_a2;
input 	input_b4;
input 	input_a3;
input 	input_b5;
input 	input_a4;
input 	input_b6;
input 	input_a5;
input 	input_b7;
input 	input_a6;
input 	input_b8;
input 	input_a7;
input 	input_b9;
input 	input_a8;
input 	input_b10;
input 	input_a9;
input 	input_b11;
input 	input_a10;
input 	input_b12;
input 	input_a11;
input 	input_b13;
input 	input_a12;
input 	input_b14;
input 	input_a13;
input 	input_b15;
input 	input_a14;
input 	input_b16;
input 	input_a15;
input 	input_b17;
input 	input_a16;
input 	input_b18;
input 	input_a17;
input 	input_b19;
input 	input_b20;
input 	input_a18;
input 	input_b21;
input 	input_a19;
input 	input_b22;
input 	input_a20;
input 	input_b23;
input 	input_a21;
input 	input_b24;
input 	input_a22;
input 	input_b25;
input 	input_a23;
input 	input_b26;
input 	input_b27;
input 	input_a24;
input 	input_b28;
input 	input_a25;
input 	input_b29;
input 	input_a26;
input 	input_b30;
input 	input_b31;
input 	input_a27;
input 	input_b32;
input 	input_b33;
input 	input_a28;
input 	input_b34;
input 	input_b35;
input 	input_a29;
input 	input_b36;
input 	input_b37;
input 	input_a30;
input 	input_b38;
input 	input_b39;
input 	input_a31;
output 	Equal0;
output 	Equal01;
output 	Equal02;
output 	Selector30;
input 	halt_reg;
output 	Selector28;
output 	Selector3;
output 	Selector22;
output 	Selector2;
output 	Selector27;
output 	Selector25;
input 	input_b40;
output 	Selector24;
output 	Selector26;
output 	Selector4;
output 	Selector16;
output 	Selector7;
output 	Selector6;
output 	Selector29;
output 	Selector15;
output 	Selector5;
output 	Selector31;
output 	Selector11;
output 	Selector10;
output 	Selector21;
output 	Selector20;
output 	Selector9;
output 	Selector8;
output 	Selector14;
output 	Selector13;
output 	Selector12;
output 	Selector23;
output 	Selector19;
output 	Selector18;
output 	Selector17;
output 	Selector0;
output 	Selector1;
output 	Equal11;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~6_combout ;
wire \Add1~20_combout ;
wire \Add1~24_combout ;
wire \Add1~26_combout ;
wire \Add1~28_combout ;
wire \Add1~32_combout ;
wire \Add1~34_combout ;
wire \Add1~36_combout ;
wire \Add0~2_combout ;
wire \ShiftLeft0~14_combout ;
wire \Selector28~4_combout ;
wire \ShiftLeft0~29_combout ;
wire \Selector3~5_combout ;
wire \Selector3~7_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \ShiftRight0~69_combout ;
wire \Selector16~6_combout ;
wire \ShiftRight0~80_combout ;
wire \Selector31~2_combout ;
wire \Selector31~3_combout ;
wire \Selector31~6_combout ;
wire \Selector21~4_combout ;
wire \Selector21~5_combout ;
wire \Selector21~6_combout ;
wire \Selector9~4_combout ;
wire \Selector13~2_combout ;
wire \Selector23~3_combout ;
wire \Selector23~4_combout ;
wire \Selector19~3_combout ;
wire \Selector19~4_combout ;
wire \Selector19~5_combout ;
wire \Selector18~1_combout ;
wire \Selector18~2_combout ;
wire \Selector17~3_combout ;
wire \Selector1~5_combout ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~0_combout ;
wire \Add0~30_combout ;
wire \Add0~32_combout ;
wire \Add0~28_combout ;
wire \Add0~24_combout ;
wire \Add0~26_combout ;
wire \Add0~22_combout ;
wire \Add0~18_combout ;
wire \Add0~20_combout ;
wire \Add0~12_combout ;
wire \Add0~14_combout ;
wire \Add0~8_combout ;
wire \Add0~6_combout ;
wire \Add0~4_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Add0~36_combout ;
wire \Add0~38_combout ;
wire \Add0~40_combout ;
wire \Add0~34_combout ;
wire \Selector0~4_combout ;
wire \Selector0~2_combout ;
wire \Selector30~2_combout ;
wire \Selector30~3_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~26_combout ;
wire \Selector22~0_combout ;
wire \ShiftRight0~27_combout ;
wire \Selector0~0_combout ;
wire \ShiftLeft0~19_combout ;
wire \ShiftLeft0~17_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~15_combout ;
wire \ShiftLeft0~16_combout ;
wire \Selector31~0_combout ;
wire \ShiftRight0~0_combout ;
wire \ShiftRight0~2_combout ;
wire \ShiftRight0~4_combout ;
wire \ShiftRight0~3_combout ;
wire \ShiftRight0~5_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~14_combout ;
wire \Selector30~0_combout ;
wire \Selector1~0_combout ;
wire \ShiftLeft0~21_combout ;
wire \Selector7~4_combout ;
wire \Selector30~1_combout ;
wire \Selector0~5_combout ;
wire \Selector30~4_combout ;
wire \Selector0~6_combout ;
wire \Add1~2_combout ;
wire \Selector0~7_combout ;
wire \Selector30~5_combout ;
wire \Selector30~6_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~23_combout ;
wire \Selector0~8_combout ;
wire \Selector28~3_combout ;
wire \Selector28~5_combout ;
wire \Selector0~10_combout ;
wire \Selector0~9_combout ;
wire \Selector28~1_combout ;
wire \Selector28~2_combout ;
wire \Selector0~14_combout ;
wire \ShiftLeft0~24_combout ;
wire \ShiftLeft0~103_combout ;
wire \Selector28~6_combout ;
wire \Selector28~7_combout ;
wire \Selector3~1_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~1_combout ;
wire \Selector28~8_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~37_combout ;
wire \Selector28~9_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~32_combout ;
wire \Selector20~0_combout ;
wire \ShiftLeft0~102_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~33_combout ;
wire \Selector15~0_combout ;
wire \Selector28~0_combout ;
wire \Selector3~0_combout ;
wire \Selector29~0_combout ;
wire \Selector0~15_combout ;
wire \Selector15~1_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~40_combout ;
wire \Selector3~2_combout ;
wire \Selector0~12_combout ;
wire \Selector0~13_combout ;
wire \Selector0~11_combout ;
wire \Selector3~3_combout ;
wire \Add1~56_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~41_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~45_combout ;
wire \ShiftLeft0~46_combout ;
wire \Selector11~2_combout ;
wire \ShiftLeft0~47_combout ;
wire \Selector3~8_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~32_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \Selector3~6_combout ;
wire \Selector3~4_combout ;
wire \Selector3~9_combout ;
wire \Selector3~10_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~51_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~48_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~53_combout ;
wire \ShiftLeft0~104_combout ;
wire \ShiftLeft0~54_combout ;
wire \Selector22~1_combout ;
wire \Selector23~0_combout ;
wire \Selector22~4_combout ;
wire \Add1~18_combout ;
wire \Selector22~5_combout ;
wire \Selector22~6_combout ;
wire \Selector15~2_combout ;
wire \Selector16~0_combout ;
wire \Selector22~2_combout ;
wire \Selector22~3_combout ;
wire \Selector22~7_combout ;
wire \Selector15~3_combout ;
wire \Selector22~8_combout ;
wire \Selector2~0_combout ;
wire \Add1~58_combout ;
wire \Selector2~1_combout ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \Selector2~6_combout ;
wire \Selector2~7_combout ;
wire \Selector27~6_combout ;
wire \Selector27~5_combout ;
wire \Selector27~7_combout ;
wire \Add1~8_combout ;
wire \Selector27~0_combout ;
wire \ShiftLeft0~40_combout ;
wire \Selector27~1_combout ;
wire \Selector7~13_combout ;
wire \Selector7~5_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~53_combout ;
wire \Selector27~2_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \Selector25~5_combout ;
wire \Selector25~4_combout ;
wire \Selector25~6_combout ;
wire \Add1~12_combout ;
wire \Selector25~0_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~73_combout ;
wire \ShiftLeft0~75_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~65_combout ;
wire \Selector25~1_combout ;
wire \Selector25~2_combout ;
wire \Selector25~3_combout ;
wire \Selector24~0_combout ;
wire \Selector0~3_combout ;
wire \Selector24~1_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \Selector24~5_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~29_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~73_combout ;
wire \Selector24~6_combout ;
wire \Selector24~7_combout ;
wire \Selector24~3_combout ;
wire \Add1~14_combout ;
wire \Selector24~2_combout ;
wire \Selector24~4_combout ;
wire \Selector26~4_combout ;
wire \Selector26~5_combout ;
wire \Selector26~6_combout ;
wire \Add1~10_combout ;
wire \Add0~10_combout ;
wire \Selector26~0_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~74_combout ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \Selector26~3_combout ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~82_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~85_combout ;
wire \Selector4~3_combout ;
wire \Selector4~4_combout ;
wire \Selector4~5_combout ;
wire \Add1~54_combout ;
wire \Selector4~6_combout ;
wire \Selector4~0_combout ;
wire \Selector16~9_combout ;
wire \Selector8~2_combout ;
wire \ShiftLeft0~88_combout ;
wire \ShiftLeft0~87_combout ;
wire \Selector16~2_combout ;
wire \Selector16~1_combout ;
wire \Selector16~3_combout ;
wire \Selector16~4_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~71_combout ;
wire \Add1~30_combout ;
wire \Selector16~5_combout ;
wire \Selector16~7_combout ;
wire \Selector16~8_combout ;
wire \Selector7~8_combout ;
wire \Selector7~6_combout ;
wire \Add1~48_combout ;
wire \Selector7~7_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~28_combout ;
wire \Selector7~9_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~78_combout ;
wire \ShiftLeft0~90_combout ;
wire \ShiftLeft0~91_combout ;
wire \Selector7~10_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~77_combout ;
wire \Selector7~11_combout ;
wire \Selector6~0_combout ;
wire \Selector6~2_combout ;
wire \ShiftLeft0~58_combout ;
wire \Selector6~3_combout ;
wire \ShiftLeft0~65_combout ;
wire \Selector6~4_combout ;
wire \Selector6~5_combout ;
wire \Add1~50_combout ;
wire \Selector6~1_combout ;
wire \Selector29~2_combout ;
wire \Selector29~3_combout ;
wire \Add1~4_combout ;
wire \Selector29~4_combout ;
wire \Selector29~5_combout ;
wire \Selector29~6_combout ;
wire \Selector29~7_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~81_combout ;
wire \Selector29~8_combout ;
wire \Selector29~9_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~68_combout ;
wire \Selector21~0_combout ;
wire \ShiftRight0~79_combout ;
wire \Selector29~1_combout ;
wire \ShiftLeft0~89_combout ;
wire \Selector15~13_combout ;
wire \Selector15~9_combout ;
wire \Selector15~11_combout ;
wire \Selector15~10_combout ;
wire \Selector15~8_combout ;
wire \Selector15~12_combout ;
wire \Selector15~4_combout ;
wire \Selector15~5_combout ;
wire \Selector15~6_combout ;
wire \Selector15~7_combout ;
wire \Selector5~0_combout ;
wire \Selector5~2_combout ;
wire \ShiftLeft0~98_combout ;
wire \ShiftLeft0~99_combout ;
wire \ShiftLeft0~100_combout ;
wire \ShiftLeft0~97_combout ;
wire \ShiftLeft0~96_combout ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \Selector5~5_combout ;
wire \Add1~52_combout ;
wire \Selector5~1_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \Selector0~16_combout ;
wire \Selector31~1_combout ;
wire \Selector31~9_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~86_combout ;
wire \Selector0~1_combout ;
wire \Selector31~4_combout ;
wire \Selector31~5_combout ;
wire \Selector31~7_combout ;
wire \Selector31~8_combout ;
wire \Selector0~17_combout ;
wire \Selector31~10_combout ;
wire \Selector11~4_combout ;
wire \Add1~40_combout ;
wire \Selector11~3_combout ;
wire \Selector11~5_combout ;
wire \Selector11~6_combout ;
wire \Selector11~10_combout ;
wire \Selector11~7_combout ;
wire \Selector11~8_combout ;
wire \Add1~42_combout ;
wire \Selector10~3_combout ;
wire \ShiftLeft0~62_combout ;
wire \ShiftLeft0~66_combout ;
wire \Selector10~4_combout ;
wire \Selector10~5_combout ;
wire \ShiftLeft0~70_combout ;
wire \Selector10~9_combout ;
wire \Selector10~6_combout ;
wire \Selector10~7_combout ;
wire \Selector21~1_combout ;
wire \Selector21~2_combout ;
wire \Selector21~3_combout ;
wire \Selector21~7_combout ;
wire \Selector21~8_combout ;
wire \Selector20~1_combout ;
wire \Selector20~4_combout ;
wire \Add1~22_combout ;
wire \Selector20~5_combout ;
wire \Selector20~6_combout ;
wire \Selector20~2_combout ;
wire \Selector20~3_combout ;
wire \Selector20~7_combout ;
wire \Selector9~0_combout ;
wire \Selector9~6_combout ;
wire \Selector9~1_combout ;
wire \Selector9~2_combout ;
wire \Add1~44_combout ;
wire \Selector9~3_combout ;
wire \Selector9~5_combout ;
wire \Selector9~7_combout ;
wire \Add1~46_combout ;
wire \Selector8~3_combout ;
wire \Selector8~4_combout ;
wire \Selector0~18_combout ;
wire \Selector8~9_combout ;
wire \Selector8~5_combout ;
wire \Selector8~6_combout ;
wire \Selector8~7_combout ;
wire \ShiftLeft0~92_combout ;
wire \Selector14~0_combout ;
wire \Selector14~1_combout ;
wire \Selector14~2_combout ;
wire \Selector14~3_combout ;
wire \Selector14~4_combout ;
wire \Selector14~5_combout ;
wire \Selector14~6_combout ;
wire \ShiftLeft0~94_combout ;
wire \ShiftLeft0~93_combout ;
wire \ShiftLeft0~95_combout ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \Selector13~4_combout ;
wire \Selector13~3_combout ;
wire \Selector13~5_combout ;
wire \Selector13~6_combout ;
wire \Selector12~0_combout ;
wire \Selector12~2_combout ;
wire \Selector12~4_combout ;
wire \Add1~38_combout ;
wire \Selector12~3_combout ;
wire \Selector12~5_combout ;
wire \Selector12~1_combout ;
wire \Selector12~6_combout ;
wire \Selector23~2_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~43_combout ;
wire \Selector23~1_combout ;
wire \Selector23~5_combout ;
wire \Add1~16_combout ;
wire \Add0~16_combout ;
wire \Selector23~6_combout ;
wire \Selector23~7_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~85_combout ;
wire \Selector23~8_combout ;
wire \Selector23~9_combout ;
wire \Selector19~7_combout ;
wire \Selector19~0_combout ;
wire \ShiftRight0~47_combout ;
wire \Selector19~1_combout ;
wire \Selector19~2_combout ;
wire \Selector19~6_combout ;
wire \Selector19~8_combout ;
wire \Selector10~2_combout ;
wire \ShiftLeft0~71_combout ;
wire \Selector18~4_combout ;
wire \Selector18~3_combout ;
wire \Selector18~5_combout ;
wire \Selector18~6_combout ;
wire \Selector18~0_combout ;
wire \Selector18~7_combout ;
wire \ShiftLeft0~101_combout ;
wire \Selector17~0_combout ;
wire \Selector17~4_combout ;
wire \Selector17~2_combout ;
wire \Selector17~5_combout ;
wire \Selector17~1_combout ;
wire \Selector17~6_combout ;
wire \Selector0~27_combout ;
wire \Selector0~20_combout ;
wire \Selector0~21_combout ;
wire \Selector1~1_combout ;
wire \ShiftLeft0~59_combout ;
wire \Selector0~22_combout ;
wire \Selector0~23_combout ;
wire \Selector0~24_combout ;
wire \Selector0~19_combout ;
wire \Selector0~25_combout ;
wire \Selector0~26_combout ;
wire \Selector1~6_combout ;
wire \Selector1~7_combout ;
wire \Selector1~3_combout ;
wire \Selector1~2_combout ;
wire \Selector1~4_combout ;
wire \Selector1~8_combout ;
wire \Selector1~9_combout ;
wire \Add1~60_combout ;
wire \Selector1~10_combout ;
wire \Equal11~10_combout ;
wire \Equal11~7_combout ;
wire \Equal11~8_combout ;
wire \Equal11~6_combout ;
wire \Equal11~9_combout ;
wire \Equal11~3_combout ;
wire \Equal11~2_combout ;
wire \Equal11~1_combout ;
wire \Equal11~4_combout ;
wire \Equal11~0_combout ;
wire \Equal11~5_combout ;


// Location: LCCOMB_X47_Y33_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\input_b~85_combout  & (\input_a~137_combout  $ (VCC))) # (!\input_b~85_combout  & ((\input_a~137_combout ) # (GND)))
// \Add1~1  = CARRY((\input_a~137_combout ) # (!\input_b~85_combout ))

	.dataa(input_b39),
	.datab(input_a31),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66DD;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\input_a~128_combout  & ((\input_b~79_combout  & (!\Add1~5 )) # (!\input_b~79_combout  & (\Add1~5  & VCC)))) # (!\input_a~128_combout  & ((\input_b~79_combout  & ((\Add1~5 ) # (GND))) # (!\input_b~79_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((\input_a~128_combout  & (\input_b~79_combout  & !\Add1~5 )) # (!\input_a~128_combout  & ((\input_b~79_combout ) # (!\Add1~5 ))))

	.dataa(input_a28),
	.datab(input_b33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h694D;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\input_b~65_combout  $ (\input_a~107_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\input_b~65_combout  & (\input_a~107_combout  & !\Add1~19 )) # (!\input_b~65_combout  & ((\input_a~107_combout ) # (!\Add1~19 ))))

	.dataa(input_b23),
	.datab(input_a21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h964D;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\input_a~101_combout  $ (\input_b~61_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\input_a~101_combout  & ((!\Add1~23 ) # (!\input_b~61_combout ))) # (!\input_a~101_combout  & (!\input_b~61_combout  & !\Add1~23 )))

	.dataa(input_a19),
	.datab(input_b21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h962B;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\input_b~59_combout  & ((\input_a~98_combout  & (!\Add1~25 )) # (!\input_a~98_combout  & ((\Add1~25 ) # (GND))))) # (!\input_b~59_combout  & ((\input_a~98_combout  & (\Add1~25  & VCC)) # (!\input_a~98_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((\input_b~59_combout  & ((!\Add1~25 ) # (!\input_a~98_combout ))) # (!\input_b~59_combout  & (!\input_a~98_combout  & !\Add1~25 )))

	.dataa(input_b20),
	.datab(input_a18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h692B;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\input_a~95_combout  $ (\input_b~57_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\input_a~95_combout  & ((!\Add1~27 ) # (!\input_b~57_combout ))) # (!\input_a~95_combout  & (!\input_b~57_combout  & !\Add1~27 )))

	.dataa(input_a17),
	.datab(input_b19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\input_b~51_combout  $ (\input_a~91_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\input_b~51_combout  & (\input_a~91_combout  & !\Add1~31 )) # (!\input_b~51_combout  & ((\input_a~91_combout ) # (!\Add1~31 ))))

	.dataa(input_b17),
	.datab(input_a15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\input_b~48_combout  & ((\input_a~89_combout  & (!\Add1~33 )) # (!\input_a~89_combout  & ((\Add1~33 ) # (GND))))) # (!\input_b~48_combout  & ((\input_a~89_combout  & (\Add1~33  & VCC)) # (!\input_a~89_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((\input_b~48_combout  & ((!\Add1~33 ) # (!\input_a~89_combout ))) # (!\input_b~48_combout  & (!\input_a~89_combout  & !\Add1~33 )))

	.dataa(input_b16),
	.datab(input_a14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h692B;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\input_b~45_combout  $ (\input_a~87_combout  $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\input_b~45_combout  & (\input_a~87_combout  & !\Add1~35 )) # (!\input_b~45_combout  & ((\input_a~87_combout ) # (!\Add1~35 ))))

	.dataa(input_b15),
	.datab(input_a13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\input_a~134_combout  & ((\input_b~83_combout  & (\Add0~1  & VCC)) # (!\input_b~83_combout  & (!\Add0~1 )))) # (!\input_a~134_combout  & ((\input_b~83_combout  & (!\Add0~1 )) # (!\input_b~83_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\input_a~134_combout  & (!\input_b~83_combout  & !\Add0~1 )) # (!\input_a~134_combout  & ((!\Add0~1 ) # (!\input_b~83_combout ))))

	.dataa(input_a30),
	.datab(input_b37),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\input_b~39_combout ) # ((\input_b~33_combout ) # ((\input_b~30_combout ) # (\input_b~36_combout )))

	.dataa(input_b13),
	.datab(input_b11),
	.datac(input_b10),
	.datad(input_b12),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N28
cycloneive_lcell_comb \Selector28~4 (
// Equation(s):
// \Selector28~4_combout  = (\Add0~6_combout  & ((\Selector0~12_combout ) # ((\Selector0~13_combout  & \Add1~6_combout )))) # (!\Add0~6_combout  & (\Selector0~13_combout  & ((\Add1~6_combout ))))

	.dataa(\Add0~6_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\Selector28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~4 .lut_mask = 16'hECA0;
defparam \Selector28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N22
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (\input_b~85_combout  & ((\input_a~69_combout ))) # (!\input_b~85_combout  & (\input_a~67_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a3),
	.datad(input_a4),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N14
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// \Selector3~5_combout  = (\Selector3~1_combout  & (((!\ShiftLeft0~103_combout )))) # (!\Selector3~1_combout  & ((\ShiftLeft0~103_combout  & (\ShiftLeft0~29_combout )) # (!\ShiftLeft0~103_combout  & ((\ShiftLeft0~28_combout )))))

	.dataa(\Selector3~1_combout ),
	.datab(\ShiftLeft0~29_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'h44FA;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N26
cycloneive_lcell_comb \Selector3~7 (
// Equation(s):
// \Selector3~7_combout  = (\input_a~67_combout  & ((\Selector0~8_combout ) # ((\input_b~15_combout  & \Selector0~9_combout )))) # (!\input_a~67_combout  & (\input_b~15_combout  & (\Selector0~8_combout )))

	.dataa(input_a3),
	.datab(input_b5),
	.datac(\Selector0~8_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~7 .lut_mask = 16'hE8E0;
defparam \Selector3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N10
cycloneive_lcell_comb \Selector2~2 (
// Equation(s):
// \Selector2~2_combout  = (\Selector3~1_combout  & (((!\ShiftLeft0~103_combout )))) # (!\Selector3~1_combout  & ((\ShiftLeft0~103_combout  & ((\ShiftLeft0~59_combout ))) # (!\ShiftLeft0~103_combout  & (\ShiftLeft0~58_combout ))))

	.dataa(\ShiftLeft0~58_combout ),
	.datab(\ShiftLeft0~59_combout ),
	.datac(\Selector3~1_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~2 .lut_mask = 16'h0CFA;
defparam \Selector2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N0
cycloneive_lcell_comb \Selector2~3 (
// Equation(s):
// \Selector2~3_combout  = (\Selector2~2_combout  & ((\ShiftLeft0~66_combout ) # ((!\Selector3~1_combout )))) # (!\Selector2~2_combout  & (((\Selector3~1_combout  & \ShiftLeft0~55_combout ))))

	.dataa(\Selector2~2_combout ),
	.datab(\ShiftLeft0~66_combout ),
	.datac(\Selector3~1_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~3 .lut_mask = 16'hDA8A;
defparam \Selector2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N0
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & (\ShiftRight0~67_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~68_combout )))))

	.dataa(\ShiftRight0~67_combout ),
	.datab(input_b33),
	.datac(input_b35),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'h2320;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \Selector16~6 (
// Equation(s):
// \Selector16~6_combout  = (\input_a~93_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_b~54_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(input_b18),
	.datad(input_a16),
	.cin(gnd),
	.combout(\Selector16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~6 .lut_mask = 16'hEA00;
defparam \Selector16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N22
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (\input_b~85_combout  & (\input_a~128_combout )) # (!\input_b~85_combout  & ((\input_a~131_combout )))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a28),
	.datad(input_a29),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N22
cycloneive_lcell_comb \Selector31~2 (
// Equation(s):
// \Selector31~2_combout  = (\Selector0~4_combout ) # (\Selector0~6_combout )

	.dataa(gnd),
	.datab(\Selector0~4_combout ),
	.datac(\Selector0~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~2 .lut_mask = 16'hFCFC;
defparam \Selector31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N16
cycloneive_lcell_comb \Selector31~3 (
// Equation(s):
// \Selector31~3_combout  = (\Add0~0_combout  & ((\Selector31~2_combout ) # ((\Selector0~7_combout  & \Add1~0_combout )))) # (!\Add0~0_combout  & (\Selector0~7_combout  & ((\Add1~0_combout ))))

	.dataa(\Add0~0_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector31~2_combout ),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\Selector31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~3 .lut_mask = 16'hECA0;
defparam \Selector31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N2
cycloneive_lcell_comb \Selector31~6 (
// Equation(s):
// \Selector31~6_combout  = (\input_b~77_combout  & ((\input_b~79_combout  & ((\ShiftRight0~77_combout ))) # (!\input_b~79_combout  & (\Selector23~1_combout ))))

	.dataa(\Selector23~1_combout ),
	.datab(input_b31),
	.datac(input_b33),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\Selector31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~6 .lut_mask = 16'hC808;
defparam \Selector31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N12
cycloneive_lcell_comb \Selector21~4 (
// Equation(s):
// \Selector21~4_combout  = (\Selector0~11_combout  & (!\input_b~65_combout  & !\input_a~107_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(input_b23),
	.datac(gnd),
	.datad(input_a21),
	.cin(gnd),
	.combout(\Selector21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~4 .lut_mask = 16'h0022;
defparam \Selector21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N26
cycloneive_lcell_comb \Selector21~5 (
// Equation(s):
// \Selector21~5_combout  = (\Add1~20_combout  & ((\Selector0~13_combout ) # ((\Add0~20_combout  & \Selector0~12_combout )))) # (!\Add1~20_combout  & (((\Add0~20_combout  & \Selector0~12_combout ))))

	.dataa(\Add1~20_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add0~20_combout ),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~5 .lut_mask = 16'hF888;
defparam \Selector21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N0
cycloneive_lcell_comb \Selector21~6 (
// Equation(s):
// \Selector21~6_combout  = (\Selector21~5_combout ) # ((\Selector21~4_combout ) # ((\Selector0~8_combout  & \input_a~107_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(input_a21),
	.datac(\Selector21~5_combout ),
	.datad(\Selector21~4_combout ),
	.cin(gnd),
	.combout(\Selector21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~6 .lut_mask = 16'hFFF8;
defparam \Selector21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N22
cycloneive_lcell_comb \Selector9~4 (
// Equation(s):
// \Selector9~4_combout  = (\Selector0~8_combout  & (((\input_a~79_combout ) # (\input_b~33_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\input_a~79_combout  & \input_b~33_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(input_a9),
	.datad(input_b11),
	.cin(gnd),
	.combout(\Selector9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~4 .lut_mask = 16'hEAA0;
defparam \Selector9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N22
cycloneive_lcell_comb \Selector13~2 (
// Equation(s):
// \Selector13~2_combout  = (\input_b~45_combout  & (!\input_a~87_combout  & ((\Selector0~10_combout )))) # (!\input_b~45_combout  & ((\input_a~87_combout  & ((\Selector0~10_combout ))) # (!\input_a~87_combout  & (\Selector0~11_combout ))))

	.dataa(input_b15),
	.datab(input_a13),
	.datac(\Selector0~11_combout ),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~2 .lut_mask = 16'h7610;
defparam \Selector13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N20
cycloneive_lcell_comb \Selector23~3 (
// Equation(s):
// \Selector23~3_combout  = (\input_b~69_combout  & ((\Selector0~8_combout ) # ((\input_a~113_combout  & \Selector0~9_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(input_a23),
	.datac(input_b25),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~3 .lut_mask = 16'hE0A0;
defparam \Selector23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N14
cycloneive_lcell_comb \Selector23~4 (
// Equation(s):
// \Selector23~4_combout  = (\Selector23~3_combout ) # ((\Selector0~10_combout  & (\input_b~69_combout  $ (\input_a~113_combout ))))

	.dataa(input_b25),
	.datab(input_a23),
	.datac(\Selector0~10_combout ),
	.datad(\Selector23~3_combout ),
	.cin(gnd),
	.combout(\Selector23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~4 .lut_mask = 16'hFF60;
defparam \Selector23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N16
cycloneive_lcell_comb \Selector19~3 (
// Equation(s):
// \Selector19~3_combout  = (!\input_b~61_combout  & (\Selector0~11_combout  & !\input_a~101_combout ))

	.dataa(gnd),
	.datab(input_b21),
	.datac(\Selector0~11_combout ),
	.datad(input_a19),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~3 .lut_mask = 16'h0030;
defparam \Selector19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N2
cycloneive_lcell_comb \Selector19~4 (
// Equation(s):
// \Selector19~4_combout  = (\Selector0~12_combout  & ((\Add0~24_combout ) # ((\Selector0~13_combout  & \Add1~24_combout )))) # (!\Selector0~12_combout  & (((\Selector0~13_combout  & \Add1~24_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~24_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Add1~24_combout ),
	.cin(gnd),
	.combout(\Selector19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~4 .lut_mask = 16'hF888;
defparam \Selector19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N12
cycloneive_lcell_comb \Selector19~5 (
// Equation(s):
// \Selector19~5_combout  = (\Selector19~3_combout ) # ((\Selector19~4_combout ) # ((\Selector0~8_combout  & \input_a~101_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector19~3_combout ),
	.datac(input_a19),
	.datad(\Selector19~4_combout ),
	.cin(gnd),
	.combout(\Selector19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~5 .lut_mask = 16'hFFEC;
defparam \Selector19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N2
cycloneive_lcell_comb \Selector18~1 (
// Equation(s):
// \Selector18~1_combout  = (\Selector0~8_combout ) # ((\input_a~98_combout  & \Selector0~9_combout ))

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(input_a18),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~1 .lut_mask = 16'hFAAA;
defparam \Selector18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \Selector18~2 (
// Equation(s):
// \Selector18~2_combout  = (\input_b~59_combout  & ((\Selector18~1_combout ) # ((!\input_a~98_combout  & \Selector0~10_combout )))) # (!\input_b~59_combout  & (((\input_a~98_combout  & \Selector0~10_combout ))))

	.dataa(input_b20),
	.datab(\Selector18~1_combout ),
	.datac(input_a18),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~2 .lut_mask = 16'hDA88;
defparam \Selector18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N10
cycloneive_lcell_comb \Selector17~3 (
// Equation(s):
// \Selector17~3_combout  = (\Selector0~12_combout  & ((\Add0~28_combout ) # ((\Selector0~13_combout  & \Add1~28_combout )))) # (!\Selector0~12_combout  & (\Selector0~13_combout  & ((\Add1~28_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add0~28_combout ),
	.datad(\Add1~28_combout ),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~3 .lut_mask = 16'hECA0;
defparam \Selector17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N8
cycloneive_lcell_comb \Selector1~5 (
// Equation(s):
// \Selector1~5_combout  = (\ShiftLeft0~104_combout  & (((\Selector1~1_combout ) # (\ShiftLeft0~29_combout )))) # (!\ShiftLeft0~104_combout  & (\input_a~63_combout  & (!\Selector1~1_combout )))

	.dataa(\ShiftLeft0~104_combout ),
	.datab(input_a1),
	.datac(\Selector1~1_combout ),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~5 .lut_mask = 16'hAEA4;
defparam \Selector1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// Add1 = \input_b~6_combout  $ (\Add1~61  $ (!\input_a~61_combout ))

	.dataa(input_b2),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(\Add1~61 ),
	.combout(Add1),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h5AA5;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// Add0 = (\input_a~81_combout  & ((\input_b~36_combout  & (\Add0~41  & VCC)) # (!\input_b~36_combout  & (!\Add0~41 )))) # (!\input_a~81_combout  & ((\input_b~36_combout  & (!\Add0~41 )) # (!\input_b~36_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\input_a~81_combout  & (!\input_b~36_combout  & !\Add0~41 )) # (!\input_a~81_combout  & ((!\Add0~41 ) # (!\input_b~36_combout ))))

	.dataa(input_a10),
	.datab(input_b12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(Add0),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// Add01 = ((\input_a~79_combout  $ (\input_b~33_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\input_a~79_combout  & ((\input_b~33_combout ) # (!\Add0~43 ))) # (!\input_a~79_combout  & (\input_b~33_combout  & !\Add0~43 )))

	.dataa(input_a9),
	.datab(input_b11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(Add01),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// Add02 = (\input_b~30_combout  & ((\input_a~77_combout  & (\Add0~45  & VCC)) # (!\input_a~77_combout  & (!\Add0~45 )))) # (!\input_b~30_combout  & ((\input_a~77_combout  & (!\Add0~45 )) # (!\input_a~77_combout  & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\input_b~30_combout  & (!\input_a~77_combout  & !\Add0~45 )) # (!\input_b~30_combout  & ((!\Add0~45 ) # (!\input_a~77_combout ))))

	.dataa(input_b10),
	.datab(input_a8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(Add02),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// Add03 = ((\input_b~27_combout  $ (\input_a~75_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\input_b~27_combout  & ((\input_a~75_combout ) # (!\Add0~47 ))) # (!\input_b~27_combout  & (\input_a~75_combout  & !\Add0~47 )))

	.dataa(input_b9),
	.datab(input_a7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(Add03),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// Add04 = (\input_b~24_combout  & ((\input_a~73_combout  & (\Add0~49  & VCC)) # (!\input_a~73_combout  & (!\Add0~49 )))) # (!\input_b~24_combout  & ((\input_a~73_combout  & (!\Add0~49 )) # (!\input_a~73_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\input_b~24_combout  & (!\input_a~73_combout  & !\Add0~49 )) # (!\input_b~24_combout  & ((!\Add0~49 ) # (!\input_a~73_combout ))))

	.dataa(input_b8),
	.datab(input_a6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(Add04),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// Add05 = ((\input_a~71_combout  $ (\input_b~21_combout  $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\input_a~71_combout  & ((\input_b~21_combout ) # (!\Add0~51 ))) # (!\input_a~71_combout  & (\input_b~21_combout  & !\Add0~51 )))

	.dataa(input_a5),
	.datab(input_b7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(Add05),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// Add06 = (\input_b~18_combout  & ((\input_a~69_combout  & (\Add0~53  & VCC)) # (!\input_a~69_combout  & (!\Add0~53 )))) # (!\input_b~18_combout  & ((\input_a~69_combout  & (!\Add0~53 )) # (!\input_a~69_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\input_b~18_combout  & (!\input_a~69_combout  & !\Add0~53 )) # (!\input_b~18_combout  & ((!\Add0~53 ) # (!\input_a~69_combout ))))

	.dataa(input_b6),
	.datab(input_a4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(Add06),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// Add07 = ((\input_b~15_combout  $ (\input_a~67_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\input_b~15_combout  & ((\input_a~67_combout ) # (!\Add0~55 ))) # (!\input_b~15_combout  & (\input_a~67_combout  & !\Add0~55 )))

	.dataa(input_b5),
	.datab(input_a3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(Add07),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// Add08 = (\input_b~12_combout  & ((\input_a~65_combout  & (\Add0~57  & VCC)) # (!\input_a~65_combout  & (!\Add0~57 )))) # (!\input_b~12_combout  & ((\input_a~65_combout  & (!\Add0~57 )) # (!\input_a~65_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\input_b~12_combout  & (!\input_a~65_combout  & !\Add0~57 )) # (!\input_b~12_combout  & ((!\Add0~57 ) # (!\input_a~65_combout ))))

	.dataa(input_b4),
	.datab(input_a2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(Add08),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// Add09 = ((\input_b~9_combout  $ (\input_a~63_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\input_b~9_combout  & ((\input_a~63_combout ) # (!\Add0~59 ))) # (!\input_b~9_combout  & (\input_a~63_combout  & !\Add0~59 )))

	.dataa(input_b3),
	.datab(input_a1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(Add09),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// Add010 = \input_b~6_combout  $ (\Add0~61  $ (\input_a~61_combout ))

	.dataa(input_b2),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(\Add0~61 ),
	.combout(Add010),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hA55A;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \out~0 (
// Equation(s):
// out = \input_a~61_combout  $ (((\input_b~5_combout ) # ((Result_EX_31 & \input_b~1_combout ))))

	.dataa(input_a),
	.datab(Result_EX_31),
	.datac(input_b),
	.datad(input_b1),
	.cin(gnd),
	.combout(out),
	.cout());
// synopsys translate_off
defparam \out~0 .lut_mask = 16'h556A;
defparam \out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N4
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// Equal0 = \input_a~61_combout  $ (\Add0~0_combout )

	.dataa(input_a),
	.datab(gnd),
	.datac(\Add0~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h5A5A;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N22
cycloneive_lcell_comb \Equal0~5 (
// Equation(s):
// Equal01 = (!\Add0~30_combout  & (!\Add0~32_combout  & (!\Add0~28_combout  & \Equal0~4_combout )))

	.dataa(\Add0~30_combout ),
	.datab(\Add0~32_combout ),
	.datac(\Add0~28_combout ),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(Equal01),
	.cout());
// synopsys translate_off
defparam \Equal0~5 .lut_mask = 16'h0100;
defparam \Equal0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N2
cycloneive_lcell_comb \Equal0~6 (
// Equation(s):
// Equal02 = (!\Add0~36_combout  & (!\Add0~38_combout  & (!\Add0~40_combout  & !\Add0~34_combout )))

	.dataa(\Add0~36_combout ),
	.datab(\Add0~38_combout ),
	.datac(\Add0~40_combout ),
	.datad(\Add0~34_combout ),
	.cin(gnd),
	.combout(Equal02),
	.cout());
// synopsys translate_off
defparam \Equal0~6 .lut_mask = 16'h0001;
defparam \Equal0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N24
cycloneive_lcell_comb \Selector30~7 (
// Equation(s):
// Selector30 = (\Selector30~3_combout ) # ((\Selector30~0_combout ) # ((\Selector30~1_combout ) # (\Selector30~6_combout )))

	.dataa(\Selector30~3_combout ),
	.datab(\Selector30~0_combout ),
	.datac(\Selector30~1_combout ),
	.datad(\Selector30~6_combout ),
	.cin(gnd),
	.combout(Selector30),
	.cout());
// synopsys translate_off
defparam \Selector30~7 .lut_mask = 16'hFFFE;
defparam \Selector30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N0
cycloneive_lcell_comb \Selector28~10 (
// Equation(s):
// Selector28 = (\Selector28~7_combout ) # ((\Selector28~0_combout ) # ((\Selector28~9_combout  & \Selector29~0_combout )))

	.dataa(\Selector28~7_combout ),
	.datab(\Selector28~9_combout ),
	.datac(\Selector28~0_combout ),
	.datad(\Selector29~0_combout ),
	.cin(gnd),
	.combout(Selector28),
	.cout());
// synopsys translate_off
defparam \Selector28~10 .lut_mask = 16'hFEFA;
defparam \Selector28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N8
cycloneive_lcell_comb \Selector3~11 (
// Equation(s):
// Selector3 = (\Selector3~2_combout ) # ((\Selector3~10_combout ) # ((Add07 & \Selector0~12_combout )))

	.dataa(Add07),
	.datab(\Selector3~2_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Selector3~10_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~11 .lut_mask = 16'hFFEC;
defparam \Selector3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N18
cycloneive_lcell_comb \Selector22~9 (
// Equation(s):
// Selector22 = (\Selector22~1_combout ) # ((\Selector22~8_combout ) # ((\ShiftRight0~20_combout  & \Selector23~0_combout )))

	.dataa(\Selector22~1_combout ),
	.datab(\ShiftRight0~20_combout ),
	.datac(\Selector23~0_combout ),
	.datad(\Selector22~8_combout ),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~9 .lut_mask = 16'hFFEA;
defparam \Selector22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N20
cycloneive_lcell_comb \Selector2~8 (
// Equation(s):
// Selector2 = (\Selector2~0_combout ) # ((\Selector2~7_combout ) # ((Add08 & \Selector0~12_combout )))

	.dataa(Add08),
	.datab(\Selector0~12_combout ),
	.datac(\Selector2~0_combout ),
	.datad(\Selector2~7_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~8 .lut_mask = 16'hFFF8;
defparam \Selector2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N0
cycloneive_lcell_comb \Selector27~8 (
// Equation(s):
// Selector27 = (\Selector27~7_combout ) # ((\Selector27~0_combout ) # (\Selector27~4_combout ))

	.dataa(\Selector27~7_combout ),
	.datab(gnd),
	.datac(\Selector27~0_combout ),
	.datad(\Selector27~4_combout ),
	.cin(gnd),
	.combout(Selector27),
	.cout());
// synopsys translate_off
defparam \Selector27~8 .lut_mask = 16'hFFFA;
defparam \Selector27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N30
cycloneive_lcell_comb \Selector25~7 (
// Equation(s):
// Selector25 = (\Selector25~6_combout ) # ((\Selector25~0_combout ) # (\Selector25~3_combout ))

	.dataa(gnd),
	.datab(\Selector25~6_combout ),
	.datac(\Selector25~0_combout ),
	.datad(\Selector25~3_combout ),
	.cin(gnd),
	.combout(Selector25),
	.cout());
// synopsys translate_off
defparam \Selector25~7 .lut_mask = 16'hFFFC;
defparam \Selector25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Selector24~8 (
// Equation(s):
// Selector24 = (\Selector24~0_combout ) # ((\Selector24~1_combout ) # ((\Selector24~7_combout ) # (\Selector24~4_combout )))

	.dataa(\Selector24~0_combout ),
	.datab(\Selector24~1_combout ),
	.datac(\Selector24~7_combout ),
	.datad(\Selector24~4_combout ),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~8 .lut_mask = 16'hFFFE;
defparam \Selector24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N14
cycloneive_lcell_comb \Selector26~7 (
// Equation(s):
// Selector26 = (\Selector26~6_combout ) # ((\Selector26~0_combout ) # (\Selector26~3_combout ))

	.dataa(\Selector26~6_combout ),
	.datab(gnd),
	.datac(\Selector26~0_combout ),
	.datad(\Selector26~3_combout ),
	.cin(gnd),
	.combout(Selector26),
	.cout());
// synopsys translate_off
defparam \Selector26~7 .lut_mask = 16'hFFFA;
defparam \Selector26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N8
cycloneive_lcell_comb \Selector4~7 (
// Equation(s):
// Selector4 = (\Selector4~6_combout ) # ((\Selector4~0_combout ) # ((Add06 & \Selector0~6_combout )))

	.dataa(Add06),
	.datab(\Selector0~6_combout ),
	.datac(\Selector4~6_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~7 .lut_mask = 16'hFFF8;
defparam \Selector4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N10
cycloneive_lcell_comb \Selector16~10 (
// Equation(s):
// Selector16 = (\Selector16~3_combout ) # ((\Selector16~8_combout ) # ((\Selector16~9_combout  & \ShiftLeft0~88_combout )))

	.dataa(\Selector16~9_combout ),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\Selector16~3_combout ),
	.datad(\Selector16~8_combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~10 .lut_mask = 16'hFFF8;
defparam \Selector16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N30
cycloneive_lcell_comb \Selector7~12 (
// Equation(s):
// Selector7 = (\Selector7~8_combout ) # ((\Selector7~6_combout ) # ((\Selector7~7_combout ) # (\Selector7~11_combout )))

	.dataa(\Selector7~8_combout ),
	.datab(\Selector7~6_combout ),
	.datac(\Selector7~7_combout ),
	.datad(\Selector7~11_combout ),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~12 .lut_mask = 16'hFFFE;
defparam \Selector7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N20
cycloneive_lcell_comb \Selector6~6 (
// Equation(s):
// Selector6 = (\Selector6~0_combout ) # ((\Selector6~2_combout ) # ((\Selector6~5_combout ) # (\Selector6~1_combout )))

	.dataa(\Selector6~0_combout ),
	.datab(\Selector6~2_combout ),
	.datac(\Selector6~5_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~6 .lut_mask = 16'hFFFE;
defparam \Selector6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N22
cycloneive_lcell_comb \Selector29~10 (
// Equation(s):
// Selector29 = (\Selector29~7_combout ) # ((\Selector29~1_combout ) # ((\Selector29~0_combout  & \Selector29~9_combout )))

	.dataa(\Selector29~7_combout ),
	.datab(\Selector29~0_combout ),
	.datac(\Selector29~9_combout ),
	.datad(\Selector29~1_combout ),
	.cin(gnd),
	.combout(Selector29),
	.cout());
// synopsys translate_off
defparam \Selector29~10 .lut_mask = 16'hFFEA;
defparam \Selector29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N28
cycloneive_lcell_comb \Selector15~14 (
// Equation(s):
// Selector15 = (\Selector15~12_combout ) # ((\Selector15~7_combout ) # ((\ShiftLeft0~89_combout  & \Selector15~13_combout )))

	.dataa(\ShiftLeft0~89_combout ),
	.datab(\Selector15~13_combout ),
	.datac(\Selector15~12_combout ),
	.datad(\Selector15~7_combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~14 .lut_mask = 16'hFFF8;
defparam \Selector15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N10
cycloneive_lcell_comb \Selector5~6 (
// Equation(s):
// Selector5 = (\Selector5~0_combout ) # ((\Selector5~2_combout ) # ((\Selector5~5_combout ) # (\Selector5~1_combout )))

	.dataa(\Selector5~0_combout ),
	.datab(\Selector5~2_combout ),
	.datac(\Selector5~5_combout ),
	.datad(\Selector5~1_combout ),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~6 .lut_mask = 16'hFFFE;
defparam \Selector5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N6
cycloneive_lcell_comb \Selector31~11 (
// Equation(s):
// Selector31 = (\Selector31~1_combout ) # ((\Selector31~10_combout ) # ((\LessThan0~62_combout  & \Selector0~16_combout )))

	.dataa(\LessThan0~62_combout ),
	.datab(\Selector0~16_combout ),
	.datac(\Selector31~1_combout ),
	.datad(\Selector31~10_combout ),
	.cin(gnd),
	.combout(Selector31),
	.cout());
// synopsys translate_off
defparam \Selector31~11 .lut_mask = 16'hFFF8;
defparam \Selector31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N18
cycloneive_lcell_comb \Selector11~9 (
// Equation(s):
// Selector11 = (\Selector11~3_combout ) # ((\Selector11~8_combout ) # ((\Selector11~4_combout  & \ShiftLeft0~40_combout )))

	.dataa(\Selector11~4_combout ),
	.datab(\ShiftLeft0~40_combout ),
	.datac(\Selector11~3_combout ),
	.datad(\Selector11~8_combout ),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~9 .lut_mask = 16'hFFF8;
defparam \Selector11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N16
cycloneive_lcell_comb \Selector10~8 (
// Equation(s):
// Selector10 = (\Selector10~3_combout ) # ((\Selector10~7_combout ) # ((\ShiftLeft0~67_combout  & \Selector11~4_combout )))

	.dataa(\ShiftLeft0~67_combout ),
	.datab(\Selector10~3_combout ),
	.datac(\Selector11~4_combout ),
	.datad(\Selector10~7_combout ),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~8 .lut_mask = 16'hFFEC;
defparam \Selector10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N10
cycloneive_lcell_comb \Selector21~9 (
// Equation(s):
// Selector21 = (\Selector21~1_combout ) # ((\Selector21~8_combout ) # ((\ShiftRight0~78_combout  & \Selector23~0_combout )))

	.dataa(\Selector21~1_combout ),
	.datab(\Selector21~8_combout ),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector23~0_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~9 .lut_mask = 16'hFEEE;
defparam \Selector21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N6
cycloneive_lcell_comb \Selector20~8 (
// Equation(s):
// Selector20 = (\Selector20~1_combout ) # ((\Selector20~7_combout ) # ((\ShiftRight0~37_combout  & \Selector16~0_combout )))

	.dataa(\ShiftRight0~37_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector20~1_combout ),
	.datad(\Selector20~7_combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
// synopsys translate_off
defparam \Selector20~8 .lut_mask = 16'hFFF8;
defparam \Selector20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N22
cycloneive_lcell_comb \Selector9~8 (
// Equation(s):
// Selector9 = (\Selector9~0_combout ) # ((\Selector9~7_combout ) # ((\ShiftLeft0~75_combout  & \Selector11~4_combout )))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(\Selector11~4_combout ),
	.datac(\Selector9~0_combout ),
	.datad(\Selector9~7_combout ),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~8 .lut_mask = 16'hFFF8;
defparam \Selector9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N20
cycloneive_lcell_comb \Selector8~8 (
// Equation(s):
// Selector8 = (\Selector8~3_combout ) # ((\Selector8~7_combout ) # ((\ShiftLeft0~77_combout  & \Selector11~4_combout )))

	.dataa(\ShiftLeft0~77_combout ),
	.datab(\Selector8~3_combout ),
	.datac(\Selector8~7_combout ),
	.datad(\Selector11~4_combout ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~8 .lut_mask = 16'hFEFC;
defparam \Selector8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N4
cycloneive_lcell_comb \Selector14~7 (
// Equation(s):
// Selector14 = (\Selector14~0_combout ) # ((\Selector14~6_combout ) # ((\ShiftLeft0~92_combout  & \Selector15~13_combout )))

	.dataa(\ShiftLeft0~92_combout ),
	.datab(\Selector14~0_combout ),
	.datac(\Selector14~6_combout ),
	.datad(\Selector15~13_combout ),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~7 .lut_mask = 16'hFEFC;
defparam \Selector14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N24
cycloneive_lcell_comb \Selector13~7 (
// Equation(s):
// Selector13 = (\Selector13~0_combout ) # ((\Selector13~6_combout ) # ((\ShiftLeft0~95_combout  & \Selector15~13_combout )))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(\Selector13~0_combout ),
	.datac(\Selector15~13_combout ),
	.datad(\Selector13~6_combout ),
	.cin(gnd),
	.combout(Selector13),
	.cout());
// synopsys translate_off
defparam \Selector13~7 .lut_mask = 16'hFFEC;
defparam \Selector13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N14
cycloneive_lcell_comb \Selector12~7 (
// Equation(s):
// Selector12 = (\Selector12~0_combout ) # ((\Selector12~6_combout ) # ((\ShiftRight0~33_combout  & \Selector15~1_combout )))

	.dataa(\Selector12~0_combout ),
	.datab(\ShiftRight0~33_combout ),
	.datac(\Selector15~1_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(Selector12),
	.cout());
// synopsys translate_off
defparam \Selector12~7 .lut_mask = 16'hFFEA;
defparam \Selector12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N30
cycloneive_lcell_comb \Selector23~10 (
// Equation(s):
// Selector23 = (\Selector23~2_combout ) # ((\Selector23~9_combout ) # ((\ShiftRight0~77_combout  & \Selector23~0_combout )))

	.dataa(\ShiftRight0~77_combout ),
	.datab(\Selector23~2_combout ),
	.datac(\Selector23~0_combout ),
	.datad(\Selector23~9_combout ),
	.cin(gnd),
	.combout(Selector23),
	.cout());
// synopsys translate_off
defparam \Selector23~10 .lut_mask = 16'hFFEC;
defparam \Selector23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N16
cycloneive_lcell_comb \Selector19~9 (
// Equation(s):
// Selector19 = (\Selector19~8_combout ) # ((\ShiftLeft0~47_combout  & \Selector16~9_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~47_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\Selector19~8_combout ),
	.cin(gnd),
	.combout(Selector19),
	.cout());
// synopsys translate_off
defparam \Selector19~9 .lut_mask = 16'hFFC0;
defparam \Selector19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N30
cycloneive_lcell_comb \Selector18~8 (
// Equation(s):
// Selector18 = (\Selector18~7_combout ) # ((\ShiftLeft0~71_combout  & \Selector16~9_combout ))

	.dataa(\ShiftLeft0~71_combout ),
	.datab(gnd),
	.datac(\Selector16~9_combout ),
	.datad(\Selector18~7_combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~8 .lut_mask = 16'hFFA0;
defparam \Selector18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N28
cycloneive_lcell_comb \Selector17~7 (
// Equation(s):
// Selector17 = (\Selector17~0_combout ) # ((\Selector17~6_combout ) # ((\ShiftLeft0~101_combout  & \Selector16~9_combout )))

	.dataa(\ShiftLeft0~101_combout ),
	.datab(\Selector17~0_combout ),
	.datac(\Selector17~6_combout ),
	.datad(\Selector16~9_combout ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~7 .lut_mask = 16'hFEFC;
defparam \Selector17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N24
cycloneive_lcell_comb \Selector0~28 (
// Equation(s):
// Selector0 = (\Selector0~27_combout ) # ((\Selector0~26_combout ) # ((\Selector0~12_combout  & Add010)))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~27_combout ),
	.datac(\Selector0~26_combout ),
	.datad(Add010),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~28 .lut_mask = 16'hFEFC;
defparam \Selector0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N14
cycloneive_lcell_comb \Selector1~11 (
// Equation(s):
// Selector1 = (\Selector1~8_combout ) # ((\Selector1~10_combout ) # ((Add09 & \Selector0~12_combout )))

	.dataa(\Selector1~8_combout ),
	.datab(Add09),
	.datac(\Selector0~12_combout ),
	.datad(\Selector1~10_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~11 .lut_mask = 16'hFFEA;
defparam \Selector1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \Equal11~11 (
// Equation(s):
// Equal11 = (!Selector31 & (\Equal11~10_combout  & (\Equal11~9_combout  & \Equal11~5_combout )))

	.dataa(Selector31),
	.datab(\Equal11~10_combout ),
	.datac(\Equal11~9_combout ),
	.datad(\Equal11~5_combout ),
	.cin(gnd),
	.combout(Equal11),
	.cout());
// synopsys translate_off
defparam \Equal11~11 .lut_mask = 16'h4000;
defparam \Equal11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\input_a~134_combout  & ((\input_b~83_combout  & (!\Add1~1 )) # (!\input_b~83_combout  & (\Add1~1  & VCC)))) # (!\input_a~134_combout  & ((\input_b~83_combout  & ((\Add1~1 ) # (GND))) # (!\input_b~83_combout  & (!\Add1~1 ))))
// \Add1~3  = CARRY((\input_a~134_combout  & (\input_b~83_combout  & !\Add1~1 )) # (!\input_a~134_combout  & ((\input_b~83_combout ) # (!\Add1~1 ))))

	.dataa(input_a30),
	.datab(input_b37),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h694D;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\input_a~131_combout  $ (\input_b~81_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\input_a~131_combout  & ((!\Add1~3 ) # (!\input_b~81_combout ))) # (!\input_a~131_combout  & (!\input_b~81_combout  & !\Add1~3 )))

	.dataa(input_a29),
	.datab(input_b35),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h962B;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\input_a~125_combout  $ (\input_b~77_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\input_a~125_combout  & ((!\Add1~7 ) # (!\input_b~77_combout ))) # (!\input_a~125_combout  & (!\input_b~77_combout  & !\Add1~7 )))

	.dataa(input_a27),
	.datab(input_b31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h962B;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\input_b~75_combout  & ((\input_a~122_combout  & (!\Add1~9 )) # (!\input_a~122_combout  & ((\Add1~9 ) # (GND))))) # (!\input_b~75_combout  & ((\input_a~122_combout  & (\Add1~9  & VCC)) # (!\input_a~122_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((\input_b~75_combout  & ((!\Add1~9 ) # (!\input_a~122_combout ))) # (!\input_b~75_combout  & (!\input_a~122_combout  & !\Add1~9 )))

	.dataa(input_b29),
	.datab(input_a26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h692B;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\input_b~73_combout  $ (\input_a~119_combout  $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\input_b~73_combout  & (\input_a~119_combout  & !\Add1~11 )) # (!\input_b~73_combout  & ((\input_a~119_combout ) # (!\Add1~11 ))))

	.dataa(input_b28),
	.datab(input_a25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h964D;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\input_b~71_combout  & ((\input_a~116_combout  & (!\Add1~13 )) # (!\input_a~116_combout  & ((\Add1~13 ) # (GND))))) # (!\input_b~71_combout  & ((\input_a~116_combout  & (\Add1~13  & VCC)) # (!\input_a~116_combout  & (!\Add1~13 ))))
// \Add1~15  = CARRY((\input_b~71_combout  & ((!\Add1~13 ) # (!\input_a~116_combout ))) # (!\input_b~71_combout  & (!\input_a~116_combout  & !\Add1~13 )))

	.dataa(input_b27),
	.datab(input_a24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h692B;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((\input_a~113_combout  $ (\input_b~69_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((\input_a~113_combout  & ((!\Add1~15 ) # (!\input_b~69_combout ))) # (!\input_a~113_combout  & (!\input_b~69_combout  & !\Add1~15 )))

	.dataa(input_a23),
	.datab(input_b25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h962B;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\input_a~110_combout  & ((\input_b~67_combout  & (!\Add1~17 )) # (!\input_b~67_combout  & (\Add1~17  & VCC)))) # (!\input_a~110_combout  & ((\input_b~67_combout  & ((\Add1~17 ) # (GND))) # (!\input_b~67_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((\input_a~110_combout  & (\input_b~67_combout  & !\Add1~17 )) # (!\input_a~110_combout  & ((\input_b~67_combout ) # (!\Add1~17 ))))

	.dataa(input_a22),
	.datab(input_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h694D;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\input_a~104_combout  & ((\input_b~63_combout  & (!\Add1~21 )) # (!\input_b~63_combout  & (\Add1~21  & VCC)))) # (!\input_a~104_combout  & ((\input_b~63_combout  & ((\Add1~21 ) # (GND))) # (!\input_b~63_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((\input_a~104_combout  & (\input_b~63_combout  & !\Add1~21 )) # (!\input_a~104_combout  & ((\input_b~63_combout ) # (!\Add1~21 ))))

	.dataa(input_a20),
	.datab(input_b22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h694D;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\input_b~54_combout  & ((\input_a~93_combout  & (!\Add1~29 )) # (!\input_a~93_combout  & ((\Add1~29 ) # (GND))))) # (!\input_b~54_combout  & ((\input_a~93_combout  & (\Add1~29  & VCC)) # (!\input_a~93_combout  & (!\Add1~29 ))))
// \Add1~31  = CARRY((\input_b~54_combout  & ((!\Add1~29 ) # (!\input_a~93_combout ))) # (!\input_b~54_combout  & (!\input_a~93_combout  & !\Add1~29 )))

	.dataa(input_b18),
	.datab(input_a16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h692B;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\input_a~85_combout  & ((\input_b~42_combout  & (!\Add1~37 )) # (!\input_b~42_combout  & (\Add1~37  & VCC)))) # (!\input_a~85_combout  & ((\input_b~42_combout  & ((\Add1~37 ) # (GND))) # (!\input_b~42_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((\input_a~85_combout  & (\input_b~42_combout  & !\Add1~37 )) # (!\input_a~85_combout  & ((\input_b~42_combout ) # (!\Add1~37 ))))

	.dataa(input_a12),
	.datab(input_b14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h694D;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\input_b~39_combout  $ (\input_a~83_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\input_b~39_combout  & (\input_a~83_combout  & !\Add1~39 )) # (!\input_b~39_combout  & ((\input_a~83_combout ) # (!\Add1~39 ))))

	.dataa(input_b13),
	.datab(input_a11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h964D;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\input_b~36_combout  & ((\input_a~81_combout  & (!\Add1~41 )) # (!\input_a~81_combout  & ((\Add1~41 ) # (GND))))) # (!\input_b~36_combout  & ((\input_a~81_combout  & (\Add1~41  & VCC)) # (!\input_a~81_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((\input_b~36_combout  & ((!\Add1~41 ) # (!\input_a~81_combout ))) # (!\input_b~36_combout  & (!\input_a~81_combout  & !\Add1~41 )))

	.dataa(input_b12),
	.datab(input_a10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h692B;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\input_a~79_combout  $ (\input_b~33_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\input_a~79_combout  & ((!\Add1~43 ) # (!\input_b~33_combout ))) # (!\input_a~79_combout  & (!\input_b~33_combout  & !\Add1~43 )))

	.dataa(input_a9),
	.datab(input_b11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h962B;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\input_a~77_combout  & ((\input_b~30_combout  & (!\Add1~45 )) # (!\input_b~30_combout  & (\Add1~45  & VCC)))) # (!\input_a~77_combout  & ((\input_b~30_combout  & ((\Add1~45 ) # (GND))) # (!\input_b~30_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((\input_a~77_combout  & (\input_b~30_combout  & !\Add1~45 )) # (!\input_a~77_combout  & ((\input_b~30_combout ) # (!\Add1~45 ))))

	.dataa(input_a8),
	.datab(input_b10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h694D;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\input_a~75_combout  $ (\input_b~27_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\input_a~75_combout  & ((!\Add1~47 ) # (!\input_b~27_combout ))) # (!\input_a~75_combout  & (!\input_b~27_combout  & !\Add1~47 )))

	.dataa(input_a7),
	.datab(input_b9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h962B;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\input_b~24_combout  & ((\input_a~73_combout  & (!\Add1~49 )) # (!\input_a~73_combout  & ((\Add1~49 ) # (GND))))) # (!\input_b~24_combout  & ((\input_a~73_combout  & (\Add1~49  & VCC)) # (!\input_a~73_combout  & (!\Add1~49 ))))
// \Add1~51  = CARRY((\input_b~24_combout  & ((!\Add1~49 ) # (!\input_a~73_combout ))) # (!\input_b~24_combout  & (!\input_a~73_combout  & !\Add1~49 )))

	.dataa(input_b8),
	.datab(input_a6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h692B;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((\input_a~71_combout  $ (\input_b~21_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((\input_a~71_combout  & ((!\Add1~51 ) # (!\input_b~21_combout ))) # (!\input_a~71_combout  & (!\input_b~21_combout  & !\Add1~51 )))

	.dataa(input_a5),
	.datab(input_b7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\input_b~18_combout  & ((\input_a~69_combout  & (!\Add1~53 )) # (!\input_a~69_combout  & ((\Add1~53 ) # (GND))))) # (!\input_b~18_combout  & ((\input_a~69_combout  & (\Add1~53  & VCC)) # (!\input_a~69_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((\input_b~18_combout  & ((!\Add1~53 ) # (!\input_a~69_combout ))) # (!\input_b~18_combout  & (!\input_a~69_combout  & !\Add1~53 )))

	.dataa(input_b6),
	.datab(input_a4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h692B;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\input_b~15_combout  $ (\input_a~67_combout  $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\input_b~15_combout  & (\input_a~67_combout  & !\Add1~55 )) # (!\input_b~15_combout  & ((\input_a~67_combout ) # (!\Add1~55 ))))

	.dataa(input_b5),
	.datab(input_a3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h964D;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (\input_a~65_combout  & ((\input_b~12_combout  & (!\Add1~57 )) # (!\input_b~12_combout  & (\Add1~57  & VCC)))) # (!\input_a~65_combout  & ((\input_b~12_combout  & ((\Add1~57 ) # (GND))) # (!\input_b~12_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((\input_a~65_combout  & (\input_b~12_combout  & !\Add1~57 )) # (!\input_a~65_combout  & ((\input_b~12_combout ) # (!\Add1~57 ))))

	.dataa(input_a2),
	.datab(input_b4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h694D;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\input_b~9_combout  $ (\input_a~63_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\input_b~9_combout  & (\input_a~63_combout  & !\Add1~59 )) # (!\input_b~9_combout  & ((\input_a~63_combout ) # (!\Add1~59 ))))

	.dataa(input_b3),
	.datab(input_a1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h964D;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\input_a~137_combout  & (\input_b~85_combout  $ (VCC))) # (!\input_a~137_combout  & (\input_b~85_combout  & VCC))
// \Add0~1  = CARRY((\input_a~137_combout  & \input_b~85_combout ))

	.dataa(input_a31),
	.datab(input_b39),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\input_a~131_combout  $ (\input_b~81_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\input_a~131_combout  & ((\input_b~81_combout ) # (!\Add0~3 ))) # (!\input_a~131_combout  & (\input_b~81_combout  & !\Add0~3 )))

	.dataa(input_a29),
	.datab(input_b35),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\input_a~128_combout  & ((\input_b~79_combout  & (\Add0~5  & VCC)) # (!\input_b~79_combout  & (!\Add0~5 )))) # (!\input_a~128_combout  & ((\input_b~79_combout  & (!\Add0~5 )) # (!\input_b~79_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\input_a~128_combout  & (!\input_b~79_combout  & !\Add0~5 )) # (!\input_a~128_combout  & ((!\Add0~5 ) # (!\input_b~79_combout ))))

	.dataa(input_a28),
	.datab(input_b33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\input_a~125_combout  $ (\input_b~77_combout  $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\input_a~125_combout  & ((\input_b~77_combout ) # (!\Add0~7 ))) # (!\input_a~125_combout  & (\input_b~77_combout  & !\Add0~7 )))

	.dataa(input_a27),
	.datab(input_b31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\input_b~75_combout  & ((\input_a~122_combout  & (\Add0~9  & VCC)) # (!\input_a~122_combout  & (!\Add0~9 )))) # (!\input_b~75_combout  & ((\input_a~122_combout  & (!\Add0~9 )) # (!\input_a~122_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\input_b~75_combout  & (!\input_a~122_combout  & !\Add0~9 )) # (!\input_b~75_combout  & ((!\Add0~9 ) # (!\input_a~122_combout ))))

	.dataa(input_b29),
	.datab(input_a26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\input_a~119_combout  $ (\input_b~73_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\input_a~119_combout  & ((\input_b~73_combout ) # (!\Add0~11 ))) # (!\input_a~119_combout  & (\input_b~73_combout  & !\Add0~11 )))

	.dataa(input_a25),
	.datab(input_b28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\input_a~116_combout  & ((\input_b~71_combout  & (\Add0~13  & VCC)) # (!\input_b~71_combout  & (!\Add0~13 )))) # (!\input_a~116_combout  & ((\input_b~71_combout  & (!\Add0~13 )) # (!\input_b~71_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\input_a~116_combout  & (!\input_b~71_combout  & !\Add0~13 )) # (!\input_a~116_combout  & ((!\Add0~13 ) # (!\input_b~71_combout ))))

	.dataa(input_a24),
	.datab(input_b27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\input_a~113_combout  $ (\input_b~69_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\input_a~113_combout  & ((\input_b~69_combout ) # (!\Add0~15 ))) # (!\input_a~113_combout  & (\input_b~69_combout  & !\Add0~15 )))

	.dataa(input_a23),
	.datab(input_b25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\input_a~110_combout  & ((\input_b~67_combout  & (\Add0~17  & VCC)) # (!\input_b~67_combout  & (!\Add0~17 )))) # (!\input_a~110_combout  & ((\input_b~67_combout  & (!\Add0~17 )) # (!\input_b~67_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\input_a~110_combout  & (!\input_b~67_combout  & !\Add0~17 )) # (!\input_a~110_combout  & ((!\Add0~17 ) # (!\input_b~67_combout ))))

	.dataa(input_a22),
	.datab(input_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\input_b~65_combout  $ (\input_a~107_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\input_b~65_combout  & ((\input_a~107_combout ) # (!\Add0~19 ))) # (!\input_b~65_combout  & (\input_a~107_combout  & !\Add0~19 )))

	.dataa(input_b23),
	.datab(input_a21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\input_b~63_combout  & ((\input_a~104_combout  & (\Add0~21  & VCC)) # (!\input_a~104_combout  & (!\Add0~21 )))) # (!\input_b~63_combout  & ((\input_a~104_combout  & (!\Add0~21 )) # (!\input_a~104_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\input_b~63_combout  & (!\input_a~104_combout  & !\Add0~21 )) # (!\input_b~63_combout  & ((!\Add0~21 ) # (!\input_a~104_combout ))))

	.dataa(input_b22),
	.datab(input_a20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\input_b~61_combout  $ (\input_a~101_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\input_b~61_combout  & ((\input_a~101_combout ) # (!\Add0~23 ))) # (!\input_b~61_combout  & (\input_a~101_combout  & !\Add0~23 )))

	.dataa(input_b21),
	.datab(input_a19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\input_b~59_combout  & ((\input_a~98_combout  & (\Add0~25  & VCC)) # (!\input_a~98_combout  & (!\Add0~25 )))) # (!\input_b~59_combout  & ((\input_a~98_combout  & (!\Add0~25 )) # (!\input_a~98_combout  & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\input_b~59_combout  & (!\input_a~98_combout  & !\Add0~25 )) # (!\input_b~59_combout  & ((!\Add0~25 ) # (!\input_a~98_combout ))))

	.dataa(input_b20),
	.datab(input_a18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\input_a~95_combout  $ (\input_b~57_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\input_a~95_combout  & ((\input_b~57_combout ) # (!\Add0~27 ))) # (!\input_a~95_combout  & (\input_b~57_combout  & !\Add0~27 )))

	.dataa(input_a17),
	.datab(input_b19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\input_b~54_combout  & ((\input_a~93_combout  & (\Add0~29  & VCC)) # (!\input_a~93_combout  & (!\Add0~29 )))) # (!\input_b~54_combout  & ((\input_a~93_combout  & (!\Add0~29 )) # (!\input_a~93_combout  & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\input_b~54_combout  & (!\input_a~93_combout  & !\Add0~29 )) # (!\input_b~54_combout  & ((!\Add0~29 ) # (!\input_a~93_combout ))))

	.dataa(input_b18),
	.datab(input_a16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\input_a~91_combout  $ (\input_b~51_combout  $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\input_a~91_combout  & ((\input_b~51_combout ) # (!\Add0~31 ))) # (!\input_a~91_combout  & (\input_b~51_combout  & !\Add0~31 )))

	.dataa(input_a15),
	.datab(input_b17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\input_a~89_combout  & ((\input_b~48_combout  & (\Add0~33  & VCC)) # (!\input_b~48_combout  & (!\Add0~33 )))) # (!\input_a~89_combout  & ((\input_b~48_combout  & (!\Add0~33 )) # (!\input_b~48_combout  & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\input_a~89_combout  & (!\input_b~48_combout  & !\Add0~33 )) # (!\input_a~89_combout  & ((!\Add0~33 ) # (!\input_b~48_combout ))))

	.dataa(input_a14),
	.datab(input_b16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\input_b~45_combout  $ (\input_a~87_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\input_b~45_combout  & ((\input_a~87_combout ) # (!\Add0~35 ))) # (!\input_b~45_combout  & (\input_a~87_combout  & !\Add0~35 )))

	.dataa(input_b15),
	.datab(input_a13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\input_b~42_combout  & ((\input_a~85_combout  & (\Add0~37  & VCC)) # (!\input_a~85_combout  & (!\Add0~37 )))) # (!\input_b~42_combout  & ((\input_a~85_combout  & (!\Add0~37 )) # (!\input_a~85_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\input_b~42_combout  & (!\input_a~85_combout  & !\Add0~37 )) # (!\input_b~42_combout  & ((!\Add0~37 ) # (!\input_a~85_combout ))))

	.dataa(input_b14),
	.datab(input_a12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\input_a~83_combout  $ (\input_b~39_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\input_a~83_combout  & ((\input_b~39_combout ) # (!\Add0~39 ))) # (!\input_a~83_combout  & (\input_b~39_combout  & !\Add0~39 )))

	.dataa(input_a11),
	.datab(input_b13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N2
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (!\Add0~2_combout  & (!\Add0~8_combout  & (!\Add0~6_combout  & !\Add0~4_combout )))

	.dataa(\Add0~2_combout ),
	.datab(\Add0~8_combout ),
	.datac(\Add0~6_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h0001;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N12
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// \Equal0~2_combout  = (!\Add0~10_combout  & (!\Add0~12_combout  & (!\Add0~14_combout  & \Equal0~1_combout )))

	.dataa(\Add0~10_combout ),
	.datab(\Add0~12_combout ),
	.datac(\Add0~14_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h0100;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N18
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// \Equal0~3_combout  = (!\Add0~16_combout  & (!\Add0~18_combout  & (!\Add0~20_combout  & \Equal0~2_combout )))

	.dataa(\Add0~16_combout ),
	.datab(\Add0~18_combout ),
	.datac(\Add0~20_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'h0100;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N28
cycloneive_lcell_comb \Equal0~4 (
// Equation(s):
// \Equal0~4_combout  = (!\Add0~24_combout  & (!\Add0~26_combout  & (!\Add0~22_combout  & \Equal0~3_combout )))

	.dataa(\Add0~24_combout ),
	.datab(\Add0~26_combout ),
	.datac(\Add0~22_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~4 .lut_mask = 16'h0100;
defparam \Equal0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N4
cycloneive_lcell_comb \Selector0~4 (
// Equation(s):
// \Selector0~4_combout  = (!ALUOP_ID_0 & (ALUOP_ID_1 & (ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~4 .lut_mask = 16'h0040;
defparam \Selector0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N16
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// \Selector0~2_combout  = (ALUOP_ID_0 & (!ALUOP_ID_1 & (ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'h0020;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N2
cycloneive_lcell_comb \Selector30~2 (
// Equation(s):
// \Selector30~2_combout  = (\Selector0~2_combout ) # ((\Selector0~3_combout  & \input_a~134_combout ))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~2_combout ),
	.datac(gnd),
	.datad(input_a30),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~2 .lut_mask = 16'hEECC;
defparam \Selector30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N16
cycloneive_lcell_comb \Selector30~3 (
// Equation(s):
// \Selector30~3_combout  = (\input_b~83_combout  & ((\Selector30~2_combout ) # ((\Selector0~4_combout  & !\input_a~134_combout )))) # (!\input_b~83_combout  & (\Selector0~4_combout  & (\input_a~134_combout )))

	.dataa(\Selector0~4_combout ),
	.datab(input_b37),
	.datac(input_a30),
	.datad(\Selector30~2_combout ),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~3 .lut_mask = 16'hEC28;
defparam \Selector30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N4
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (\input_b~85_combout  & (\input_a~67_combout )) # (!\input_b~85_combout  & ((\input_a~69_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a3),
	.datad(input_a4),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N28
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\input_b~83_combout  & ((\ShiftRight0~17_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~18_combout ))

	.dataa(\ShiftRight0~18_combout ),
	.datab(input_b37),
	.datac(\ShiftRight0~17_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hE2E2;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N16
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (!\input_b~85_combout  & ((\input_b~83_combout  & (\input_a~61_combout )) # (!\input_b~83_combout  & ((\input_a~65_combout )))))

	.dataa(input_a),
	.datab(input_b37),
	.datac(input_a2),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'h00B8;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N18
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (\ShiftRight0~15_combout ) # ((\input_a~63_combout  & (!\input_b~83_combout  & \input_b~85_combout )))

	.dataa(input_a1),
	.datab(\ShiftRight0~15_combout ),
	.datac(input_b37),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'hCECC;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N2
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (\input_b~81_combout  & ((\ShiftRight0~16_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~19_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~19_combout ),
	.datac(input_b35),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N20
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (\input_b~85_combout  & ((\input_a~75_combout ))) # (!\input_b~85_combout  & (\input_a~77_combout ))

	.dataa(input_a8),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a7),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hEE22;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N26
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (\input_b~83_combout  & ((\ShiftRight0~21_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~22_combout ))

	.dataa(\ShiftRight0~22_combout ),
	.datab(\ShiftRight0~21_combout ),
	.datac(input_b37),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hCACA;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N30
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\input_b~85_combout  & ((\input_a~87_combout ))) # (!\input_b~85_combout  & (\input_a~89_combout ))

	.dataa(input_a14),
	.datab(input_a13),
	.datac(gnd),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hCCAA;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N12
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\input_b~85_combout  & ((\input_a~83_combout ))) # (!\input_b~85_combout  & (\input_a~85_combout ))

	.dataa(input_a12),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a11),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hEE22;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N16
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\input_b~83_combout  & ((\ShiftRight0~24_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~25_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~25_combout ),
	.datac(input_b37),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N0
cycloneive_lcell_comb \Selector22~0 (
// Equation(s):
// \Selector22~0_combout  = (\input_b~81_combout  & (\ShiftRight0~23_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~26_combout )))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftRight0~23_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~0 .lut_mask = 16'hF3C0;
defparam \Selector22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N12
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (\input_b~79_combout  & (\ShiftRight0~20_combout )) # (!\input_b~79_combout  & ((\Selector22~0_combout )))

	.dataa(input_b33),
	.datab(\ShiftRight0~20_combout ),
	.datac(\Selector22~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hD8D8;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N24
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = (!ALUOP_ID_2 & (!ALUOP_ID_1 & (ALUOP_ID_0 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_0),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'h0010;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\input_b~73_combout ) # ((\input_b~71_combout ) # (\input_b~75_combout ))

	.dataa(input_b28),
	.datab(gnd),
	.datac(input_b27),
	.datad(input_b29),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hFFFA;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N14
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\input_b~59_combout ) # ((\input_b~61_combout ) # ((\input_b~57_combout ) # (\input_b~54_combout )))

	.dataa(input_b20),
	.datab(input_b21),
	.datac(input_b19),
	.datad(input_b18),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N28
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\input_b~63_combout ) # ((\input_b~67_combout ) # ((\input_b~69_combout ) # (\input_b~65_combout )))

	.dataa(input_b22),
	.datab(input_b24),
	.datac(input_b25),
	.datad(input_b23),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N4
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (\ShiftLeft0~19_combout ) # ((\ShiftLeft0~17_combout ) # (\ShiftLeft0~18_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~19_combout ),
	.datac(\ShiftLeft0~17_combout ),
	.datad(\ShiftLeft0~18_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'hFFFC;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N30
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\input_b~27_combout ) # ((\input_b~24_combout ) # ((\input_b~18_combout ) # (\input_b~21_combout )))

	.dataa(input_b9),
	.datab(input_b8),
	.datac(input_b6),
	.datad(input_b7),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N16
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\input_b~12_combout ) # ((\input_b~15_combout ) # ((\input_b~9_combout ) # (\input_b~6_combout )))

	.dataa(input_b4),
	.datab(input_b5),
	.datac(input_b3),
	.datad(input_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N4
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (\input_b~45_combout ) # ((\input_b~42_combout ) # ((\input_b~48_combout ) # (\input_b~51_combout )))

	.dataa(input_b15),
	.datab(input_b14),
	.datac(input_b16),
	.datad(input_b17),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N12
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (\ShiftLeft0~14_combout ) # ((\ShiftLeft0~13_combout ) # ((\ShiftLeft0~12_combout ) # (\ShiftLeft0~15_combout )))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(\ShiftLeft0~13_combout ),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N2
cycloneive_lcell_comb \Selector31~0 (
// Equation(s):
// \Selector31~0_combout  = (\Selector0~0_combout  & (!\ShiftLeft0~20_combout  & !\ShiftLeft0~16_combout ))

	.dataa(gnd),
	.datab(\Selector0~0_combout ),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~0 .lut_mask = 16'h000C;
defparam \Selector31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N24
cycloneive_lcell_comb \ShiftRight0~0 (
// Equation(s):
// \ShiftRight0~0_combout  = (!\input_b~83_combout  & ((\input_b~85_combout  & (\input_a~131_combout )) # (!\input_b~85_combout  & ((\input_a~134_combout )))))

	.dataa(input_b37),
	.datab(input_a29),
	.datac(input_a30),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~0_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~0 .lut_mask = 16'h4450;
defparam \ShiftRight0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N8
cycloneive_lcell_comb \ShiftRight0~2 (
// Equation(s):
// \ShiftRight0~2_combout  = (!\input_b~81_combout  & ((\ShiftRight0~0_combout ) # ((\ShiftRight0~1_combout  & \input_b~83_combout ))))

	.dataa(\ShiftRight0~1_combout ),
	.datab(input_b37),
	.datac(input_b35),
	.datad(\ShiftRight0~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~2 .lut_mask = 16'h0F08;
defparam \ShiftRight0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N14
cycloneive_lcell_comb \ShiftRight0~4 (
// Equation(s):
// \ShiftRight0~4_combout  = (\input_b~85_combout  & ((\input_a~119_combout ))) # (!\input_b~85_combout  & (\input_a~122_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a26),
	.datad(input_a25),
	.cin(gnd),
	.combout(\ShiftRight0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~4 .lut_mask = 16'hFC30;
defparam \ShiftRight0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N24
cycloneive_lcell_comb \ShiftRight0~3 (
// Equation(s):
// \ShiftRight0~3_combout  = (\input_b~85_combout  & (\input_a~113_combout )) # (!\input_b~85_combout  & ((\input_a~116_combout )))

	.dataa(gnd),
	.datab(input_a23),
	.datac(input_a24),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~3 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N8
cycloneive_lcell_comb \ShiftRight0~5 (
// Equation(s):
// \ShiftRight0~5_combout  = (\input_b~83_combout  & ((\ShiftRight0~3_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~4_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~4_combout ),
	.datad(\ShiftRight0~3_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~5 .lut_mask = 16'hFA50;
defparam \ShiftRight0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N28
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (!\input_b~79_combout  & ((\ShiftRight0~2_combout ) # ((\input_b~81_combout  & \ShiftRight0~5_combout ))))

	.dataa(input_b33),
	.datab(input_b35),
	.datac(\ShiftRight0~2_combout ),
	.datad(\ShiftRight0~5_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'h5450;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N26
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (\input_b~85_combout  & ((\input_a~95_combout ))) # (!\input_b~85_combout  & (\input_a~98_combout ))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a18),
	.datad(input_a17),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'hFA50;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N12
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\input_b~85_combout  & (\input_a~91_combout )) # (!\input_b~85_combout  & ((\input_a~93_combout )))

	.dataa(input_b39),
	.datab(input_a15),
	.datac(input_a16),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hD8D8;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N16
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\input_b~83_combout  & ((\ShiftRight0~7_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~8_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~8_combout ),
	.datad(\ShiftRight0~7_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hFA50;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N4
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\input_b~85_combout  & ((\input_a~101_combout ))) # (!\input_b~85_combout  & (\input_a~104_combout ))

	.dataa(gnd),
	.datab(input_a20),
	.datac(input_a19),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N16
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (\input_b~83_combout  & ((\ShiftRight0~10_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~11_combout ))

	.dataa(\ShiftRight0~11_combout ),
	.datab(input_b37),
	.datac(\ShiftRight0~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'hE2E2;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N22
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\input_b~81_combout  & (\ShiftRight0~9_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~12_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~9_combout ),
	.datac(\ShiftRight0~12_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N10
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (!\input_b~77_combout  & ((\ShiftRight0~6_combout ) # ((\input_b~79_combout  & \ShiftRight0~13_combout ))))

	.dataa(input_b31),
	.datab(\ShiftRight0~6_combout ),
	.datac(input_b33),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'h5444;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N16
cycloneive_lcell_comb \Selector30~0 (
// Equation(s):
// \Selector30~0_combout  = (\Selector31~0_combout  & ((\ShiftRight0~14_combout ) # ((\ShiftRight0~27_combout  & \input_b~77_combout ))))

	.dataa(\ShiftRight0~27_combout ),
	.datab(input_b31),
	.datac(\Selector31~0_combout ),
	.datad(\ShiftRight0~14_combout ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~0 .lut_mask = 16'hF080;
defparam \Selector30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N14
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (!\input_b~83_combout  & (!\input_b~81_combout  & !\input_b~79_combout ))

	.dataa(gnd),
	.datab(input_b37),
	.datac(input_b35),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'h0003;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N4
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (\input_b~85_combout  & (\input_a~137_combout )) # (!\input_b~85_combout  & ((\input_a~134_combout )))

	.dataa(input_a31),
	.datab(gnd),
	.datac(input_b39),
	.datad(input_a30),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N8
cycloneive_lcell_comb \Selector7~4 (
// Equation(s):
// \Selector7~4_combout  = (\Selector0~1_combout  & (!\ShiftLeft0~20_combout  & !\ShiftLeft0~16_combout ))

	.dataa(\Selector0~1_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~4 .lut_mask = 16'h000A;
defparam \Selector7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N14
cycloneive_lcell_comb \Selector30~1 (
// Equation(s):
// \Selector30~1_combout  = (\Selector1~0_combout  & (\ShiftLeft0~21_combout  & (\Selector7~4_combout  & !\input_b~77_combout )))

	.dataa(\Selector1~0_combout ),
	.datab(\ShiftLeft0~21_combout ),
	.datac(\Selector7~4_combout ),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~1 .lut_mask = 16'h0080;
defparam \Selector30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N18
cycloneive_lcell_comb \Selector0~5 (
// Equation(s):
// \Selector0~5_combout  = (ALUOP_ID_0 & (ALUOP_ID_1 & (ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~5 .lut_mask = 16'h0080;
defparam \Selector0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N26
cycloneive_lcell_comb \Selector30~4 (
// Equation(s):
// \Selector30~4_combout  = (!\input_a~134_combout  & (\Selector0~5_combout  & !\input_b~83_combout ))

	.dataa(input_a30),
	.datab(\Selector0~5_combout ),
	.datac(gnd),
	.datad(input_b37),
	.cin(gnd),
	.combout(\Selector30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~4 .lut_mask = 16'h0044;
defparam \Selector30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N0
cycloneive_lcell_comb \Selector0~6 (
// Equation(s):
// \Selector0~6_combout  = (!ALUOP_ID_2 & (!ALUOP_ID_0 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~6 .lut_mask = 16'h0010;
defparam \Selector0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N10
cycloneive_lcell_comb \Selector0~7 (
// Equation(s):
// \Selector0~7_combout  = (!ALUOP_ID_2 & (ALUOP_ID_0 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~7 .lut_mask = 16'h0040;
defparam \Selector0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N28
cycloneive_lcell_comb \Selector30~5 (
// Equation(s):
// \Selector30~5_combout  = (\Add0~2_combout  & ((\Selector0~6_combout ) # ((\Add1~2_combout  & \Selector0~7_combout )))) # (!\Add0~2_combout  & (((\Add1~2_combout  & \Selector0~7_combout ))))

	.dataa(\Add0~2_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~2_combout ),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~5 .lut_mask = 16'hF888;
defparam \Selector30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N12
cycloneive_lcell_comb \Selector30~6 (
// Equation(s):
// \Selector30~6_combout  = (\Selector30~4_combout ) # ((\Selector30~5_combout ) # ((\input_a~134_combout  & \Selector0~2_combout )))

	.dataa(\Selector30~4_combout ),
	.datab(input_a30),
	.datac(\Selector0~2_combout ),
	.datad(\Selector30~5_combout ),
	.cin(gnd),
	.combout(\Selector30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~6 .lut_mask = 16'hFFEA;
defparam \Selector30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N0
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (\input_b~85_combout  & ((\input_a~131_combout ))) # (!\input_b~85_combout  & (\input_a~128_combout ))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a28),
	.datad(input_a29),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\input_b~83_combout  & (\ShiftLeft0~21_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~22_combout )))

	.dataa(input_b37),
	.datab(\ShiftLeft0~21_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N20
cycloneive_lcell_comb \Selector0~8 (
// Equation(s):
// \Selector0~8_combout  = (ALUOP_ID_2 & (ALUOP_ID_0 & (!ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~8 .lut_mask = 16'h0008;
defparam \Selector0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N20
cycloneive_lcell_comb \Selector28~3 (
// Equation(s):
// \Selector28~3_combout  = (\Selector0~11_combout  & (!\input_a~128_combout  & !\input_b~79_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(gnd),
	.datac(input_a28),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~3 .lut_mask = 16'h000A;
defparam \Selector28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N14
cycloneive_lcell_comb \Selector28~5 (
// Equation(s):
// \Selector28~5_combout  = (\Selector28~4_combout ) # ((\Selector28~3_combout ) # ((\Selector0~8_combout  & \input_a~128_combout )))

	.dataa(\Selector28~4_combout ),
	.datab(\Selector0~8_combout ),
	.datac(input_a28),
	.datad(\Selector28~3_combout ),
	.cin(gnd),
	.combout(\Selector28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~5 .lut_mask = 16'hFFEA;
defparam \Selector28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N16
cycloneive_lcell_comb \Selector0~10 (
// Equation(s):
// \Selector0~10_combout  = (ALUOP_ID_2 & (!ALUOP_ID_0 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~10 .lut_mask = 16'h0020;
defparam \Selector0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N30
cycloneive_lcell_comb \Selector0~9 (
// Equation(s):
// \Selector0~9_combout  = (ALUOP_ID_2 & (!ALUOP_ID_0 & (!ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~9 .lut_mask = 16'h0002;
defparam \Selector0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N12
cycloneive_lcell_comb \Selector28~1 (
// Equation(s):
// \Selector28~1_combout  = (\Selector0~8_combout ) # ((\input_a~128_combout  & \Selector0~9_combout ))

	.dataa(input_a28),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~1 .lut_mask = 16'hECEC;
defparam \Selector28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N26
cycloneive_lcell_comb \Selector28~2 (
// Equation(s):
// \Selector28~2_combout  = (\input_b~79_combout  & ((\Selector28~1_combout ) # ((!\input_a~128_combout  & \Selector0~10_combout )))) # (!\input_b~79_combout  & (\input_a~128_combout  & (\Selector0~10_combout )))

	.dataa(input_a28),
	.datab(input_b33),
	.datac(\Selector0~10_combout ),
	.datad(\Selector28~1_combout ),
	.cin(gnd),
	.combout(\Selector28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~2 .lut_mask = 16'hEC60;
defparam \Selector28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N30
cycloneive_lcell_comb \Selector0~14 (
// Equation(s):
// \Selector0~14_combout  = (!ALUOP_ID_0 & (!ALUOP_ID_1 & (!ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~14 .lut_mask = 16'h0001;
defparam \Selector0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N22
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (\ShiftLeft0~17_combout ) # ((\ShiftLeft0~18_combout ) # ((\ShiftLeft0~19_combout ) # (\ShiftLeft0~16_combout )))

	.dataa(\ShiftLeft0~17_combout ),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N6
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (!\input_b~78_combout  & (!\input_b~81_combout  & ((!\input_b~1_combout ) # (!Result_EX_3))))

	.dataa(input_b32),
	.datab(Result_EX_3),
	.datac(input_b),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'h0015;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N6
cycloneive_lcell_comb \Selector28~6 (
// Equation(s):
// \Selector28~6_combout  = (!\input_b~77_combout  & (\Selector0~14_combout  & (!\ShiftLeft0~24_combout  & \ShiftLeft0~103_combout )))

	.dataa(input_b31),
	.datab(\Selector0~14_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~6 .lut_mask = 16'h0400;
defparam \Selector28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N24
cycloneive_lcell_comb \Selector28~7 (
// Equation(s):
// \Selector28~7_combout  = (\Selector28~5_combout ) # ((\Selector28~2_combout ) # ((\ShiftLeft0~23_combout  & \Selector28~6_combout )))

	.dataa(\ShiftLeft0~23_combout ),
	.datab(\Selector28~5_combout ),
	.datac(\Selector28~2_combout ),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~7 .lut_mask = 16'hFEFC;
defparam \Selector28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N6
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (\input_b~79_combout ) # ((!\input_b~81_combout  & \input_b~83_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(input_b37),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'hFF30;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N10
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\input_b~85_combout  & (\input_a~107_combout )) # (!\input_b~85_combout  & ((\input_a~110_combout )))

	.dataa(input_a21),
	.datab(gnd),
	.datac(input_a22),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N18
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\input_b~83_combout  & (\ShiftRight0~11_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~3_combout )))

	.dataa(input_b37),
	.datab(\ShiftRight0~11_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~3_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hDD88;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N22
cycloneive_lcell_comb \ShiftRight0~1 (
// Equation(s):
// \ShiftRight0~1_combout  = (\input_b~85_combout  & ((\input_a~125_combout ))) # (!\input_b~85_combout  & (\input_a~128_combout ))

	.dataa(input_a28),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a27),
	.cin(gnd),
	.combout(\ShiftRight0~1_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~1 .lut_mask = 16'hEE22;
defparam \ShiftRight0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N0
cycloneive_lcell_comb \Selector28~8 (
// Equation(s):
// \Selector28~8_combout  = (\Selector3~1_combout  & (((!\ShiftLeft0~103_combout )))) # (!\Selector3~1_combout  & ((\ShiftLeft0~103_combout  & ((\ShiftRight0~1_combout ))) # (!\ShiftLeft0~103_combout  & (\ShiftRight0~34_combout ))))

	.dataa(\Selector3~1_combout ),
	.datab(\ShiftRight0~34_combout ),
	.datac(\ShiftRight0~1_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~8 .lut_mask = 16'h50EE;
defparam \Selector28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N2
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (\input_b~83_combout  & (\ShiftRight0~8_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~10_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~8_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N2
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (\input_b~81_combout  & (\ShiftRight0~35_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~36_combout )))

	.dataa(\ShiftRight0~35_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~36_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N20
cycloneive_lcell_comb \Selector28~9 (
// Equation(s):
// \Selector28~9_combout  = (\Selector3~1_combout  & ((\Selector28~8_combout  & ((\ShiftRight0~37_combout ))) # (!\Selector28~8_combout  & (\ShiftRight0~4_combout )))) # (!\Selector3~1_combout  & (\Selector28~8_combout ))

	.dataa(\Selector3~1_combout ),
	.datab(\Selector28~8_combout ),
	.datac(\ShiftRight0~4_combout ),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\Selector28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~9 .lut_mask = 16'hEC64;
defparam \Selector28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N22
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\input_b~85_combout  & (\input_a~71_combout )) # (!\input_b~85_combout  & ((\input_a~73_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a5),
	.datad(input_a6),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N24
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\input_b~83_combout  & (\ShiftRight0~18_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~21_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~18_combout ),
	.datad(\ShiftRight0~21_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N0
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\input_b~85_combout  & (\input_a~79_combout )) # (!\input_b~85_combout  & ((\input_a~81_combout )))

	.dataa(input_a9),
	.datab(gnd),
	.datac(input_a10),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N20
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (\input_b~83_combout  & (\ShiftRight0~22_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~24_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~22_combout ),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N26
cycloneive_lcell_comb \Selector20~0 (
// Equation(s):
// \Selector20~0_combout  = (\input_b~81_combout  & (\ShiftRight0~31_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~32_combout )))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftRight0~31_combout ),
	.datad(\ShiftRight0~32_combout ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~0 .lut_mask = 16'hF3C0;
defparam \Selector20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N30
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (!\input_b~82_combout  & (!\input_b~85_combout  & ((!\input_b~1_combout ) # (!Result_EX_1))))

	.dataa(Result_EX_1),
	.datab(input_b36),
	.datac(input_b39),
	.datad(input_b),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'h0103;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N0
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (\input_b~81_combout  & (((\input_a~61_combout  & \ShiftLeft0~102_combout )))) # (!\input_b~81_combout  & (\ShiftRight0~29_combout ))

	.dataa(\ShiftRight0~29_combout ),
	.datab(input_b35),
	.datac(input_a),
	.datad(\ShiftLeft0~102_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'hE222;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N12
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\input_b~79_combout  & ((\ShiftRight0~30_combout ))) # (!\input_b~79_combout  & (\Selector20~0_combout ))

	.dataa(input_b33),
	.datab(gnd),
	.datac(\Selector20~0_combout ),
	.datad(\ShiftRight0~30_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hFA50;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N28
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// \Selector15~0_combout  = (\halt_reg~10_combout  & (!ALUOP_ID_1 & (!\ShiftLeft0~20_combout  & !\ShiftLeft0~16_combout )))

	.dataa(halt_reg),
	.datab(ALUOP_ID_1),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'h0002;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N14
cycloneive_lcell_comb \Selector28~0 (
// Equation(s):
// \Selector28~0_combout  = (\ShiftRight0~33_combout  & (ALUOP_ID_0 & (\input_b~77_combout  & \Selector15~0_combout )))

	.dataa(\ShiftRight0~33_combout ),
	.datab(ALUOP_ID_0),
	.datac(input_b31),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~0 .lut_mask = 16'h8000;
defparam \Selector28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N0
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (ALUOP_ID_1) # ((ALUOP_ID_2) # ((!\ShiftLeft0~24_combout  & \input_b~77_combout )))

	.dataa(ALUOP_ID_1),
	.datab(ALUOP_ID_2),
	.datac(\ShiftLeft0~24_combout ),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hEFEE;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N22
cycloneive_lcell_comb \Selector29~0 (
// Equation(s):
// \Selector29~0_combout  = (!\ShiftLeft0~24_combout  & (!ALUOP_ID_3 & (ALUOP_ID_0 & !\Selector3~0_combout )))

	.dataa(\ShiftLeft0~24_combout ),
	.datab(ALUOP_ID_3),
	.datac(ALUOP_ID_0),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~0 .lut_mask = 16'h0010;
defparam \Selector29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N16
cycloneive_lcell_comb \Selector0~15 (
// Equation(s):
// \Selector0~15_combout  = (!ALUOP_ID_2 & (!ALUOP_ID_1 & (ALUOP_ID_0 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_0),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~15 .lut_mask = 16'h0010;
defparam \Selector0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N26
cycloneive_lcell_comb \Selector15~1 (
// Equation(s):
// \Selector15~1_combout  = (!\ShiftLeft0~16_combout  & (\Selector0~15_combout  & (!\ShiftLeft0~20_combout  & !\input_b~77_combout )))

	.dataa(\ShiftLeft0~16_combout ),
	.datab(\Selector0~15_combout ),
	.datac(\ShiftLeft0~20_combout ),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~1 .lut_mask = 16'h0004;
defparam \Selector15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N4
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\input_b~85_combout  & (\input_a~61_combout )) # (!\input_b~85_combout  & ((\input_a~63_combout )))

	.dataa(input_a),
	.datab(input_b39),
	.datac(input_a1),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hB8B8;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N28
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\input_b~85_combout  & ((\input_a~65_combout ))) # (!\input_b~85_combout  & (\input_a~67_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a3),
	.datad(input_a2),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hFC30;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N22
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\input_b~83_combout  & (\ShiftRight0~38_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~39_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~38_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N14
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\Selector15~1_combout  & (\ShiftLeft0~103_combout  & \ShiftRight0~40_combout ))

	.dataa(\Selector15~1_combout ),
	.datab(\ShiftLeft0~103_combout ),
	.datac(\ShiftRight0~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'h8080;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N28
cycloneive_lcell_comb \Selector0~12 (
// Equation(s):
// \Selector0~12_combout  = (!ALUOP_ID_0 & (ALUOP_ID_1 & (!ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~12 .lut_mask = 16'h0004;
defparam \Selector0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N24
cycloneive_lcell_comb \Selector0~13 (
// Equation(s):
// \Selector0~13_combout  = (!ALUOP_ID_2 & (ALUOP_ID_0 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~13 .lut_mask = 16'h0040;
defparam \Selector0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N22
cycloneive_lcell_comb \Selector0~11 (
// Equation(s):
// \Selector0~11_combout  = (ALUOP_ID_2 & (ALUOP_ID_0 & (ALUOP_ID_1 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~11 .lut_mask = 16'h0080;
defparam \Selector0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N24
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\input_a~67_combout  & (((!\input_b~15_combout  & \Selector0~10_combout )))) # (!\input_a~67_combout  & ((\input_b~15_combout  & ((\Selector0~10_combout ))) # (!\input_b~15_combout  & (\Selector0~11_combout ))))

	.dataa(input_a3),
	.datab(\Selector0~11_combout ),
	.datac(input_b5),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'h5E04;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N24
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\input_b~85_combout  & (\input_a~116_combout )) # (!\input_b~85_combout  & ((\input_a~113_combout )))

	.dataa(input_a24),
	.datab(gnd),
	.datac(input_a23),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N18
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\input_b~85_combout  & ((\input_a~122_combout ))) # (!\input_b~85_combout  & (\input_a~119_combout ))

	.dataa(input_a25),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a26),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hEE22;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N16
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\input_b~83_combout  & ((\ShiftLeft0~41_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~42_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~42_combout ),
	.datac(input_b37),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N30
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\input_b~85_combout  & ((\input_a~110_combout ))) # (!\input_b~85_combout  & (\input_a~107_combout ))

	.dataa(input_a21),
	.datab(gnd),
	.datac(input_a22),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N20
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\input_b~85_combout  & ((\input_a~104_combout ))) # (!\input_b~85_combout  & (\input_a~101_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a19),
	.datad(input_a20),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N2
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\input_b~83_combout  & (\ShiftLeft0~44_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~45_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N24
cycloneive_lcell_comb \Selector11~2 (
// Equation(s):
// \Selector11~2_combout  = (\input_b~81_combout  & (\ShiftLeft0~43_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~46_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~2 .lut_mask = 16'hF5A0;
defparam \Selector11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N22
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\input_b~79_combout  & (\ShiftLeft0~40_combout )) # (!\input_b~79_combout  & ((\Selector11~2_combout )))

	.dataa(\ShiftLeft0~40_combout ),
	.datab(input_b33),
	.datac(gnd),
	.datad(\Selector11~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N24
cycloneive_lcell_comb \Selector3~8 (
// Equation(s):
// \Selector3~8_combout  = (!ALUOP_ID_0 & (\input_b~77_combout  & (\ShiftLeft0~47_combout  & \Selector15~0_combout )))

	.dataa(ALUOP_ID_0),
	.datab(input_b31),
	.datac(\ShiftLeft0~47_combout ),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~8 .lut_mask = 16'h4000;
defparam \Selector3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N4
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\input_b~85_combout  & ((\input_a~73_combout ))) # (!\input_b~85_combout  & (\input_a~71_combout ))

	.dataa(input_b39),
	.datab(input_a5),
	.datac(gnd),
	.datad(input_a6),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N10
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (\input_b~85_combout  & (\input_a~93_combout )) # (!\input_b~85_combout  & ((\input_a~91_combout )))

	.dataa(gnd),
	.datab(input_a16),
	.datac(input_b39),
	.datad(input_a15),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N0
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\input_b~85_combout  & (\input_a~98_combout )) # (!\input_b~85_combout  & ((\input_a~95_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a18),
	.datad(input_a17),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N14
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\input_b~83_combout  & ((\ShiftLeft0~30_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~31_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N20
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\input_b~85_combout  & ((\input_a~85_combout ))) # (!\input_b~85_combout  & (\input_a~83_combout ))

	.dataa(gnd),
	.datab(input_a11),
	.datac(input_b39),
	.datad(input_a12),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N24
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (\input_b~85_combout  & (\input_a~89_combout )) # (!\input_b~85_combout  & ((\input_a~87_combout )))

	.dataa(input_a14),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a13),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N24
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\input_b~83_combout  & ((\ShiftLeft0~33_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~34_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N22
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (\input_b~81_combout  & (\ShiftLeft0~32_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~35_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N26
cycloneive_lcell_comb \Selector3~6 (
// Equation(s):
// \Selector3~6_combout  = (\Selector3~5_combout  & (((\ShiftLeft0~36_combout ) # (!\Selector3~1_combout )))) # (!\Selector3~5_combout  & (\ShiftLeft0~25_combout  & (\Selector3~1_combout )))

	.dataa(\Selector3~5_combout ),
	.datab(\ShiftLeft0~25_combout ),
	.datac(\Selector3~1_combout ),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~6 .lut_mask = 16'hEA4A;
defparam \Selector3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N20
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (!ALUOP_ID_0 & (!ALUOP_ID_3 & (!\ShiftLeft0~24_combout  & !\Selector3~0_combout )))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_3),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'h0001;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N16
cycloneive_lcell_comb \Selector3~9 (
// Equation(s):
// \Selector3~9_combout  = (\Selector3~7_combout ) # ((\Selector3~8_combout ) # ((\Selector3~6_combout  & \Selector3~4_combout )))

	.dataa(\Selector3~7_combout ),
	.datab(\Selector3~8_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\Selector3~4_combout ),
	.cin(gnd),
	.combout(\Selector3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~9 .lut_mask = 16'hFEEE;
defparam \Selector3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N6
cycloneive_lcell_comb \Selector3~10 (
// Equation(s):
// \Selector3~10_combout  = (\Selector3~3_combout ) # ((\Selector3~9_combout ) # ((\Selector0~13_combout  & \Add1~56_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector3~3_combout ),
	.datac(\Add1~56_combout ),
	.datad(\Selector3~9_combout ),
	.cin(gnd),
	.combout(\Selector3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~10 .lut_mask = 16'hFFEC;
defparam \Selector3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N26
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (\input_b~85_combout  & ((\input_a~119_combout ))) # (!\input_b~85_combout  & (\input_a~116_combout ))

	.dataa(input_a24),
	.datab(gnd),
	.datac(input_a25),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N12
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\input_b~85_combout  & ((\input_a~113_combout ))) # (!\input_b~85_combout  & (\input_a~110_combout ))

	.dataa(gnd),
	.datab(input_a22),
	.datac(input_a23),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N30
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\input_b~83_combout  & (\ShiftLeft0~50_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~51_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftLeft0~50_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N8
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\input_b~85_combout  & (\input_a~125_combout )) # (!\input_b~85_combout  & ((\input_a~122_combout )))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a27),
	.datad(input_a26),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N30
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\input_b~83_combout  & ((\ShiftLeft0~22_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~48_combout ))

	.dataa(input_b37),
	.datab(\ShiftLeft0~48_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N8
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & ((\ShiftLeft0~49_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~52_combout ))))

	.dataa(input_b33),
	.datab(input_b35),
	.datac(\ShiftLeft0~52_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'h5410;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N4
cycloneive_lcell_comb \ShiftLeft0~104 (
// Equation(s):
// \ShiftLeft0~104_combout  = (\input_b~80_combout ) # ((\input_b~83_combout ) # ((Result_EX_2 & \input_b~1_combout )))

	.dataa(input_b34),
	.datab(Result_EX_2),
	.datac(input_b37),
	.datad(input_b),
	.cin(gnd),
	.combout(\ShiftLeft0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~104 .lut_mask = 16'hFEFA;
defparam \ShiftLeft0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N10
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\ShiftLeft0~53_combout ) # ((\input_b~79_combout  & (\ShiftLeft0~21_combout  & !\ShiftLeft0~104_combout )))

	.dataa(input_b33),
	.datab(\ShiftLeft0~21_combout ),
	.datac(\ShiftLeft0~53_combout ),
	.datad(\ShiftLeft0~104_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hF0F8;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N4
cycloneive_lcell_comb \Selector22~1 (
// Equation(s):
// \Selector22~1_combout  = (!\input_b~77_combout  & (\Selector0~14_combout  & (!\ShiftLeft0~24_combout  & \ShiftLeft0~54_combout )))

	.dataa(input_b31),
	.datab(\Selector0~14_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~1 .lut_mask = 16'h0400;
defparam \Selector22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N8
cycloneive_lcell_comb \Selector23~0 (
// Equation(s):
// \Selector23~0_combout  = (!\input_b~79_combout  & (ALUOP_ID_0 & (\input_b~77_combout  & \Selector15~0_combout )))

	.dataa(input_b33),
	.datab(ALUOP_ID_0),
	.datac(input_b31),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~0 .lut_mask = 16'h4000;
defparam \Selector23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N18
cycloneive_lcell_comb \Selector22~4 (
// Equation(s):
// \Selector22~4_combout  = (!\input_b~67_combout  & (!\input_a~110_combout  & \Selector0~11_combout ))

	.dataa(gnd),
	.datab(input_b24),
	.datac(input_a22),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~4 .lut_mask = 16'h0300;
defparam \Selector22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N24
cycloneive_lcell_comb \Selector22~5 (
// Equation(s):
// \Selector22~5_combout  = (\Selector0~13_combout  & ((\Add1~18_combout ) # ((\Selector0~12_combout  & \Add0~18_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & (\Add0~18_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~18_combout ),
	.datad(\Add1~18_combout ),
	.cin(gnd),
	.combout(\Selector22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~5 .lut_mask = 16'hEAC0;
defparam \Selector22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N14
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// \Selector22~6_combout  = (\Selector22~4_combout ) # ((\Selector22~5_combout ) # ((\Selector0~8_combout  & \input_a~110_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector22~4_combout ),
	.datac(input_a22),
	.datad(\Selector22~5_combout ),
	.cin(gnd),
	.combout(\Selector22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hFFEC;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N20
cycloneive_lcell_comb \Selector15~2 (
// Equation(s):
// \Selector15~2_combout  = (ALUOP_ID_1) # ((!\ShiftLeft0~24_combout  & ((\input_b~79_combout ) # (\input_b~77_combout ))))

	.dataa(input_b33),
	.datab(ALUOP_ID_1),
	.datac(\ShiftLeft0~24_combout ),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~2 .lut_mask = 16'hCFCE;
defparam \Selector15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N18
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// \Selector16~0_combout  = (\halt_reg~10_combout  & (ALUOP_ID_0 & (!\ShiftLeft0~24_combout  & !\Selector15~2_combout )))

	.dataa(halt_reg),
	.datab(ALUOP_ID_0),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\Selector15~2_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'h0008;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N26
cycloneive_lcell_comb \Selector22~2 (
// Equation(s):
// \Selector22~2_combout  = (\Selector0~8_combout ) # ((\input_a~110_combout  & \Selector0~9_combout ))

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(input_a22),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~2 .lut_mask = 16'hFAAA;
defparam \Selector22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N8
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (\input_b~67_combout  & ((\Selector22~2_combout ) # ((!\input_a~110_combout  & \Selector0~10_combout )))) # (!\input_b~67_combout  & (\input_a~110_combout  & (\Selector0~10_combout )))

	.dataa(input_a22),
	.datab(\Selector0~10_combout ),
	.datac(\Selector22~2_combout ),
	.datad(input_b24),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'hF488;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N20
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// \Selector22~7_combout  = (\Selector22~6_combout ) # ((\Selector22~3_combout ) # ((\ShiftRight0~13_combout  & \Selector16~0_combout )))

	.dataa(\ShiftRight0~13_combout ),
	.datab(\Selector22~6_combout ),
	.datac(\Selector16~0_combout ),
	.datad(\Selector22~3_combout ),
	.cin(gnd),
	.combout(\Selector22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hFFEC;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N16
cycloneive_lcell_comb \Selector15~3 (
// Equation(s):
// \Selector15~3_combout  = (\input_b~79_combout  & (ALUOP_ID_0 & (!\input_b~77_combout  & \Selector15~0_combout )))

	.dataa(input_b33),
	.datab(ALUOP_ID_0),
	.datac(input_b31),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~3 .lut_mask = 16'h0800;
defparam \Selector15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N6
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// \Selector22~8_combout  = (\Selector22~7_combout ) # ((\Selector22~0_combout  & \Selector15~3_combout ))

	.dataa(\Selector22~0_combout ),
	.datab(gnd),
	.datac(\Selector22~7_combout ),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'hFAF0;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N26
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// \Selector2~0_combout  = (\ShiftRight0~16_combout  & (\ShiftLeft0~103_combout  & \Selector15~1_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~16_combout ),
	.datac(\ShiftLeft0~103_combout ),
	.datad(\Selector15~1_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'hC000;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N14
cycloneive_lcell_comb \Selector2~1 (
// Equation(s):
// \Selector2~1_combout  = (\input_b~12_combout  & (\Selector0~10_combout  & ((!\input_a~65_combout )))) # (!\input_b~12_combout  & ((\input_a~65_combout  & (\Selector0~10_combout )) # (!\input_a~65_combout  & ((\Selector0~11_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~11_combout ),
	.datac(input_b4),
	.datad(input_a2),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~1 .lut_mask = 16'h0AAC;
defparam \Selector2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N20
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// \Selector2~4_combout  = (\input_b~12_combout  & ((\Selector0~8_combout ) # ((\input_a~65_combout  & \Selector0~9_combout )))) # (!\input_b~12_combout  & (\input_a~65_combout  & (\Selector0~8_combout )))

	.dataa(input_b4),
	.datab(input_a2),
	.datac(\Selector0~8_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'hE8E0;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N0
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// \Selector2~5_combout  = (\ShiftLeft0~71_combout  & (\input_b~77_combout  & (!ALUOP_ID_0 & \Selector15~0_combout )))

	.dataa(\ShiftLeft0~71_combout ),
	.datab(input_b31),
	.datac(ALUOP_ID_0),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'h0800;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N2
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (\Selector2~4_combout ) # ((\Selector2~5_combout ) # ((\Selector2~3_combout  & \Selector3~4_combout )))

	.dataa(\Selector2~3_combout ),
	.datab(\Selector2~4_combout ),
	.datac(\Selector2~5_combout ),
	.datad(\Selector3~4_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'hFEFC;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N12
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\Selector2~1_combout ) # ((\Selector2~6_combout ) # ((\Selector0~13_combout  & \Add1~58_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Add1~58_combout ),
	.datac(\Selector2~1_combout ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'hFFF8;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N30
cycloneive_lcell_comb \Selector27~6 (
// Equation(s):
// \Selector27~6_combout  = (\input_b~77_combout  & ((\Selector0~2_combout ) # (!\input_a~125_combout ))) # (!\input_b~77_combout  & ((\input_a~125_combout )))

	.dataa(input_b31),
	.datab(\Selector0~2_combout ),
	.datac(gnd),
	.datad(input_a27),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~6 .lut_mask = 16'hDDAA;
defparam \Selector27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N20
cycloneive_lcell_comb \Selector27~5 (
// Equation(s):
// \Selector27~5_combout  = (\input_a~125_combout  & (\Selector0~3_combout )) # (!\input_a~125_combout  & ((\Selector0~5_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(gnd),
	.datac(\Selector0~5_combout ),
	.datad(input_a27),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~5 .lut_mask = 16'hAAF0;
defparam \Selector27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N8
cycloneive_lcell_comb \Selector27~7 (
// Equation(s):
// \Selector27~7_combout  = (\Selector27~6_combout  & ((\Selector0~4_combout ) # ((\Selector0~2_combout )))) # (!\Selector27~6_combout  & (((\Selector27~5_combout ))))

	.dataa(\Selector27~6_combout ),
	.datab(\Selector0~4_combout ),
	.datac(\Selector0~2_combout ),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(\Selector27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~7 .lut_mask = 16'hFDA8;
defparam \Selector27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N14
cycloneive_lcell_comb \Selector27~0 (
// Equation(s):
// \Selector27~0_combout  = (\Add0~8_combout  & ((\Selector0~6_combout ) # ((\Add1~8_combout  & \Selector0~7_combout )))) # (!\Add0~8_combout  & (((\Add1~8_combout  & \Selector0~7_combout ))))

	.dataa(\Add0~8_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~8_combout ),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~0 .lut_mask = 16'hF888;
defparam \Selector27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\input_b~81_combout  & (((\ShiftLeft0~102_combout  & \input_a~137_combout )))) # (!\input_b~81_combout  & (\ShiftLeft0~39_combout ))

	.dataa(\ShiftLeft0~39_combout ),
	.datab(input_b35),
	.datac(\ShiftLeft0~102_combout ),
	.datad(input_a31),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hE222;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N0
cycloneive_lcell_comb \Selector27~1 (
// Equation(s):
// \Selector27~1_combout  = (\Selector0~1_combout  & (!\input_b~77_combout  & (!\ShiftLeft0~24_combout  & !\input_b~79_combout )))

	.dataa(\Selector0~1_combout ),
	.datab(input_b31),
	.datac(\ShiftLeft0~24_combout ),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~1 .lut_mask = 16'h0002;
defparam \Selector27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N14
cycloneive_lcell_comb \Selector7~13 (
// Equation(s):
// \Selector7~13_combout  = (\input_b~76_combout ) # ((\input_b~79_combout ) # ((\input_b~1_combout  & Result_EX_4)))

	.dataa(input_b),
	.datab(input_b30),
	.datac(Result_EX_4),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~13 .lut_mask = 16'hFFEC;
defparam \Selector7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N4
cycloneive_lcell_comb \Selector7~5 (
// Equation(s):
// \Selector7~5_combout  = (\input_b~77_combout ) # ((\input_b~81_combout  & !\input_b~79_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(input_b33),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~5 .lut_mask = 16'hFF0C;
defparam \Selector7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N0
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\input_b~85_combout  & ((\input_a~116_combout ))) # (!\input_b~85_combout  & (\input_a~119_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a25),
	.datad(input_a24),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hFC30;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N20
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\input_b~85_combout  & (\input_a~122_combout )) # (!\input_b~85_combout  & ((\input_a~125_combout )))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a26),
	.datad(input_a27),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N22
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\input_b~83_combout  & (\ShiftRight0~51_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~52_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N26
cycloneive_lcell_comb \Selector27~2 (
// Equation(s):
// \Selector27~2_combout  = (\Selector7~5_combout  & ((\ShiftRight0~50_combout ) # ((\Selector7~13_combout )))) # (!\Selector7~5_combout  & (((\ShiftRight0~53_combout  & !\Selector7~13_combout ))))

	.dataa(\ShiftRight0~50_combout ),
	.datab(\Selector7~5_combout ),
	.datac(\ShiftRight0~53_combout ),
	.datad(\Selector7~13_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~2 .lut_mask = 16'hCCB8;
defparam \Selector27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N4
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\input_b~85_combout  & ((\input_a~77_combout ))) # (!\input_b~85_combout  & (\input_a~79_combout ))

	.dataa(input_a9),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a8),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hEE22;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N14
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\input_b~85_combout  & (\input_a~81_combout )) # (!\input_b~85_combout  & ((\input_a~83_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a10),
	.datad(input_a11),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N8
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\input_b~83_combout  & (\ShiftRight0~57_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~58_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~57_combout ),
	.datac(\ShiftRight0~58_combout ),
	.datad(input_b37),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N2
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & (\ShiftRight0~56_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~59_combout )))))

	.dataa(\ShiftRight0~56_combout ),
	.datab(input_b35),
	.datac(input_b33),
	.datad(\ShiftRight0~59_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'h0B08;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N8
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (\ShiftRight0~60_combout ) # ((\input_b~79_combout  & (\ShiftRight0~40_combout  & !\input_b~81_combout )))

	.dataa(input_b33),
	.datab(\ShiftRight0~60_combout ),
	.datac(\ShiftRight0~40_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hCCEC;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N8
cycloneive_lcell_comb \Selector27~3 (
// Equation(s):
// \Selector27~3_combout  = (\Selector7~13_combout  & ((\Selector27~2_combout  & ((\ShiftRight0~61_combout ))) # (!\Selector27~2_combout  & (\ShiftRight0~47_combout )))) # (!\Selector7~13_combout  & (((\Selector27~2_combout ))))

	.dataa(\ShiftRight0~47_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\Selector27~2_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~3 .lut_mask = 16'hF838;
defparam \Selector27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N2
cycloneive_lcell_comb \Selector27~4 (
// Equation(s):
// \Selector27~4_combout  = (\ShiftLeft0~40_combout  & ((\Selector27~1_combout ) # ((\Selector27~3_combout  & \Selector31~0_combout )))) # (!\ShiftLeft0~40_combout  & (((\Selector27~3_combout  & \Selector31~0_combout ))))

	.dataa(\ShiftLeft0~40_combout ),
	.datab(\Selector27~1_combout ),
	.datac(\Selector27~3_combout ),
	.datad(\Selector31~0_combout ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~4 .lut_mask = 16'hF888;
defparam \Selector27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N12
cycloneive_lcell_comb \Selector25~5 (
// Equation(s):
// \Selector25~5_combout  = (\input_a~119_combout  & ((\Selector0~2_combout ) # (!\input_b~73_combout ))) # (!\input_a~119_combout  & ((\input_b~73_combout )))

	.dataa(input_a25),
	.datab(\Selector0~2_combout ),
	.datac(gnd),
	.datad(input_b28),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~5 .lut_mask = 16'hDDAA;
defparam \Selector25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N14
cycloneive_lcell_comb \Selector25~4 (
// Equation(s):
// \Selector25~4_combout  = (\input_a~119_combout  & (\Selector0~3_combout )) # (!\input_a~119_combout  & ((\Selector0~5_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~5_combout ),
	.datac(input_a25),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~4 .lut_mask = 16'hACAC;
defparam \Selector25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N26
cycloneive_lcell_comb \Selector25~6 (
// Equation(s):
// \Selector25~6_combout  = (\Selector25~5_combout  & ((\Selector0~4_combout ) # ((\Selector0~2_combout )))) # (!\Selector25~5_combout  & (((\Selector25~4_combout ))))

	.dataa(\Selector25~5_combout ),
	.datab(\Selector0~4_combout ),
	.datac(\Selector25~4_combout ),
	.datad(\Selector0~2_combout ),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~6 .lut_mask = 16'hFAD8;
defparam \Selector25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N20
cycloneive_lcell_comb \Selector25~0 (
// Equation(s):
// \Selector25~0_combout  = (\Add0~12_combout  & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add1~12_combout )))) # (!\Add0~12_combout  & (\Selector0~7_combout  & ((\Add1~12_combout ))))

	.dataa(\Add0~12_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~0 .lut_mask = 16'hECA0;
defparam \Selector25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N0
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\input_b~85_combout  & (\input_a~128_combout )) # (!\input_b~85_combout  & ((\input_a~125_combout )))

	.dataa(input_a28),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a27),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N6
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\input_b~83_combout  & ((\ShiftLeft0~38_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~41_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~41_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N14
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (!\input_b~85_combout  & ((\input_b~83_combout  & (\input_a~137_combout )) # (!\input_b~83_combout  & ((\input_a~131_combout )))))

	.dataa(input_b37),
	.datab(input_b39),
	.datac(input_a31),
	.datad(input_a29),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'h3120;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N4
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\ShiftLeft0~72_combout ) # ((!\input_b~83_combout  & (\input_a~134_combout  & \input_b~85_combout )))

	.dataa(input_b37),
	.datab(input_a30),
	.datac(\ShiftLeft0~72_combout ),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hF4F0;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N12
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\input_b~81_combout  & ((\ShiftLeft0~73_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~74_combout ))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N16
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\ShiftRight0~69_combout ) # ((\ShiftRight0~38_combout  & (!\ShiftLeft0~104_combout  & \input_b~79_combout )))

	.dataa(\ShiftRight0~69_combout ),
	.datab(\ShiftRight0~38_combout ),
	.datac(\ShiftLeft0~104_combout ),
	.datad(input_b33),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hAEAA;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N8
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\input_b~85_combout  & ((\input_a~110_combout ))) # (!\input_b~85_combout  & (\input_a~113_combout ))

	.dataa(gnd),
	.datab(input_a23),
	.datac(input_a22),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N0
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\input_b~83_combout  & ((\ShiftRight0~49_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~51_combout ))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hFC30;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N6
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\input_b~83_combout  & ((\ShiftRight0~58_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~41_combout ))

	.dataa(\ShiftRight0~41_combout ),
	.datab(input_b37),
	.datac(gnd),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hEE22;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N14
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (\input_b~85_combout  & ((\input_a~89_combout ))) # (!\input_b~85_combout  & (\input_a~91_combout ))

	.dataa(gnd),
	.datab(input_a15),
	.datac(input_a14),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N28
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (\input_b~85_combout  & (\input_a~93_combout )) # (!\input_b~85_combout  & ((\input_a~95_combout )))

	.dataa(input_a16),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a17),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'hBB88;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N4
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (\input_b~83_combout  & (\ShiftRight0~42_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~44_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~42_combout ),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N0
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\input_b~81_combout  & (\ShiftRight0~63_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~64_combout )))

	.dataa(input_b35),
	.datab(\ShiftRight0~63_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~64_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hDD88;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N14
cycloneive_lcell_comb \Selector25~1 (
// Equation(s):
// \Selector25~1_combout  = (\Selector7~5_combout  & (((\Selector7~13_combout )))) # (!\Selector7~5_combout  & ((\Selector7~13_combout  & ((\ShiftRight0~65_combout ))) # (!\Selector7~13_combout  & (\ShiftRight0~66_combout ))))

	.dataa(\Selector7~5_combout ),
	.datab(\ShiftRight0~66_combout ),
	.datac(\Selector7~13_combout ),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~1 .lut_mask = 16'hF4A4;
defparam \Selector25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N18
cycloneive_lcell_comb \Selector25~2 (
// Equation(s):
// \Selector25~2_combout  = (\Selector25~1_combout  & (((\ShiftRight0~70_combout ) # (!\Selector7~5_combout )))) # (!\Selector25~1_combout  & (\ShiftRight0~62_combout  & ((\Selector7~5_combout ))))

	.dataa(\ShiftRight0~62_combout ),
	.datab(\ShiftRight0~70_combout ),
	.datac(\Selector25~1_combout ),
	.datad(\Selector7~5_combout ),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~2 .lut_mask = 16'hCAF0;
defparam \Selector25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N6
cycloneive_lcell_comb \Selector25~3 (
// Equation(s):
// \Selector25~3_combout  = (\Selector27~1_combout  & ((\ShiftLeft0~75_combout ) # ((\Selector31~0_combout  & \Selector25~2_combout )))) # (!\Selector27~1_combout  & (((\Selector31~0_combout  & \Selector25~2_combout ))))

	.dataa(\Selector27~1_combout ),
	.datab(\ShiftLeft0~75_combout ),
	.datac(\Selector31~0_combout ),
	.datad(\Selector25~2_combout ),
	.cin(gnd),
	.combout(\Selector25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~3 .lut_mask = 16'hF888;
defparam \Selector25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// \Selector24~0_combout  = (\Selector0~4_combout  & (\input_a~116_combout  $ (((\input_b~70_combout ) # (\input_b~86_combout )))))

	.dataa(\Selector0~4_combout ),
	.datab(input_a24),
	.datac(input_b26),
	.datad(input_b40),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h2228;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N10
cycloneive_lcell_comb \Selector0~3 (
// Equation(s):
// \Selector0~3_combout  = (!ALUOP_ID_0 & (!ALUOP_ID_1 & (ALUOP_ID_2 & !ALUOP_ID_3)))

	.dataa(ALUOP_ID_0),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_2),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~3 .lut_mask = 16'h0010;
defparam \Selector0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \Selector24~1 (
// Equation(s):
// \Selector24~1_combout  = (\input_b~71_combout  & ((\Selector0~2_combout ) # ((\input_a~116_combout  & \Selector0~3_combout ))))

	.dataa(input_b27),
	.datab(input_a24),
	.datac(\Selector0~2_combout ),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~1 .lut_mask = 16'hA8A0;
defparam \Selector24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N14
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\input_b~83_combout  & ((\ShiftLeft0~48_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~50_combout ))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftLeft0~50_combout ),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N2
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\input_b~81_combout  & (\ShiftLeft0~23_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~76_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N4
cycloneive_lcell_comb \Selector24~5 (
// Equation(s):
// \Selector24~5_combout  = (\Selector7~5_combout  & ((\Selector7~13_combout ) # ((\ShiftRight0~36_combout )))) # (!\Selector7~5_combout  & (!\Selector7~13_combout  & ((\ShiftRight0~34_combout ))))

	.dataa(\Selector7~5_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\ShiftRight0~36_combout ),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\Selector24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~5 .lut_mask = 16'hB9A8;
defparam \Selector24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N0
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\input_b~83_combout  & ((\input_b~85_combout  & ((\input_a~63_combout ))) # (!\input_b~85_combout  & (\input_a~65_combout ))))

	.dataa(input_a2),
	.datab(input_b37),
	.datac(input_a1),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hC088;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N10
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\ShiftRight0~28_combout ) # ((!\input_b~83_combout  & \ShiftRight0~17_combout ))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~17_combout ),
	.datad(\ShiftRight0~28_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hFF30;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N12
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\ShiftLeft0~78_combout  & ((\input_a~61_combout ) # ((\ShiftLeft0~103_combout  & \ShiftRight0~31_combout )))) # (!\ShiftLeft0~78_combout  & (\ShiftLeft0~103_combout  & ((\ShiftRight0~31_combout ))))

	.dataa(\ShiftLeft0~78_combout ),
	.datab(\ShiftLeft0~103_combout ),
	.datac(input_a),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hECA0;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N6
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (\ShiftRight0~72_combout ) # ((\input_b~81_combout  & (!\input_b~79_combout  & \ShiftRight0~29_combout )))

	.dataa(input_b35),
	.datab(input_b33),
	.datac(\ShiftRight0~29_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hFF20;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N16
cycloneive_lcell_comb \Selector24~6 (
// Equation(s):
// \Selector24~6_combout  = (\Selector7~13_combout  & ((\Selector24~5_combout  & ((\ShiftRight0~73_combout ))) # (!\Selector24~5_combout  & (\ShiftRight0~71_combout )))) # (!\Selector7~13_combout  & (((\Selector24~5_combout ))))

	.dataa(\ShiftRight0~71_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\Selector24~5_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\Selector24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~6 .lut_mask = 16'hF838;
defparam \Selector24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N6
cycloneive_lcell_comb \Selector24~7 (
// Equation(s):
// \Selector24~7_combout  = (\Selector31~0_combout  & ((\Selector24~6_combout ) # ((\ShiftLeft0~77_combout  & \Selector27~1_combout )))) # (!\Selector31~0_combout  & (\ShiftLeft0~77_combout  & ((\Selector27~1_combout ))))

	.dataa(\Selector31~0_combout ),
	.datab(\ShiftLeft0~77_combout ),
	.datac(\Selector24~6_combout ),
	.datad(\Selector27~1_combout ),
	.cin(gnd),
	.combout(\Selector24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~7 .lut_mask = 16'hECA0;
defparam \Selector24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Selector24~3 (
// Equation(s):
// \Selector24~3_combout  = (!\input_b~70_combout  & (\Selector0~5_combout  & ((!Result_EX_7) # (!\input_b~1_combout ))))

	.dataa(input_b26),
	.datab(\Selector0~5_combout ),
	.datac(input_b),
	.datad(Result_EX_7),
	.cin(gnd),
	.combout(\Selector24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~3 .lut_mask = 16'h0444;
defparam \Selector24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N22
cycloneive_lcell_comb \Selector24~2 (
// Equation(s):
// \Selector24~2_combout  = (\Selector0~7_combout  & ((\Add1~14_combout ) # ((\Selector0~6_combout  & \Add0~14_combout )))) # (!\Selector0~7_combout  & (\Selector0~6_combout  & ((\Add0~14_combout ))))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~14_combout ),
	.datad(\Add0~14_combout ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~2 .lut_mask = 16'hECA0;
defparam \Selector24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \Selector24~4 (
// Equation(s):
// \Selector24~4_combout  = (\Selector24~2_combout ) # ((\input_a~116_combout  & ((\Selector0~2_combout ))) # (!\input_a~116_combout  & (\Selector24~3_combout )))

	.dataa(\Selector24~3_combout ),
	.datab(input_a24),
	.datac(\Selector0~2_combout ),
	.datad(\Selector24~2_combout ),
	.cin(gnd),
	.combout(\Selector24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~4 .lut_mask = 16'hFFE2;
defparam \Selector24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \Selector26~4 (
// Equation(s):
// \Selector26~4_combout  = (\input_a~122_combout  & (\Selector0~3_combout )) # (!\input_a~122_combout  & ((\Selector0~5_combout )))

	.dataa(gnd),
	.datab(input_a26),
	.datac(\Selector0~3_combout ),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~4 .lut_mask = 16'hF3C0;
defparam \Selector26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Selector26~5 (
// Equation(s):
// \Selector26~5_combout  = (\input_b~75_combout  & ((\Selector0~2_combout ) # (!\input_a~122_combout ))) # (!\input_b~75_combout  & ((\input_a~122_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(input_b29),
	.datac(gnd),
	.datad(input_a26),
	.cin(gnd),
	.combout(\Selector26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~5 .lut_mask = 16'hBBCC;
defparam \Selector26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \Selector26~6 (
// Equation(s):
// \Selector26~6_combout  = (\Selector26~5_combout  & (((\Selector0~2_combout ) # (\Selector0~4_combout )))) # (!\Selector26~5_combout  & (\Selector26~4_combout ))

	.dataa(\Selector26~4_combout ),
	.datab(\Selector0~2_combout ),
	.datac(\Selector26~5_combout ),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~6 .lut_mask = 16'hFACA;
defparam \Selector26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N6
cycloneive_lcell_comb \Selector26~0 (
// Equation(s):
// \Selector26~0_combout  = (\Add1~10_combout  & ((\Selector0~7_combout ) # ((\Selector0~6_combout  & \Add0~10_combout )))) # (!\Add1~10_combout  & (((\Selector0~6_combout  & \Add0~10_combout ))))

	.dataa(\Add1~10_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~0 .lut_mask = 16'hF888;
defparam \Selector26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N4
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\input_b~81_combout  & (!\input_b~83_combout  & (\ShiftLeft0~21_combout ))) # (!\input_b~81_combout  & (((\ShiftLeft0~49_combout ))))

	.dataa(input_b37),
	.datab(\ShiftLeft0~21_combout ),
	.datac(\ShiftLeft0~49_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'h44F0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N8
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & ((\ShiftRight0~19_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~23_combout ))))

	.dataa(input_b33),
	.datab(input_b35),
	.datac(\ShiftRight0~23_combout ),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'h5410;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y29_N30
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\ShiftRight0~75_combout ) # ((\input_b~79_combout  & (!\input_b~81_combout  & \ShiftRight0~16_combout )))

	.dataa(input_b33),
	.datab(input_b35),
	.datac(\ShiftRight0~75_combout ),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hF2F0;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N4
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (\input_b~81_combout  & ((\ShiftRight0~26_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~9_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftRight0~9_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hFC30;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N16
cycloneive_lcell_comb \Selector26~1 (
// Equation(s):
// \Selector26~1_combout  = (\Selector7~13_combout  & (((\Selector7~5_combout ) # (\ShiftRight0~74_combout )))) # (!\Selector7~13_combout  & (\ShiftRight0~5_combout  & (!\Selector7~5_combout )))

	.dataa(\ShiftRight0~5_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\Selector7~5_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~1 .lut_mask = 16'hCEC2;
defparam \Selector26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N18
cycloneive_lcell_comb \Selector26~2 (
// Equation(s):
// \Selector26~2_combout  = (\Selector7~5_combout  & ((\Selector26~1_combout  & ((\ShiftRight0~76_combout ))) # (!\Selector26~1_combout  & (\ShiftRight0~12_combout )))) # (!\Selector7~5_combout  & (((\Selector26~1_combout ))))

	.dataa(\ShiftRight0~12_combout ),
	.datab(\Selector7~5_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\Selector26~1_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~2 .lut_mask = 16'hF388;
defparam \Selector26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N24
cycloneive_lcell_comb \Selector26~3 (
// Equation(s):
// \Selector26~3_combout  = (\Selector31~0_combout  & ((\Selector26~2_combout ) # ((\Selector27~1_combout  & \ShiftLeft0~67_combout )))) # (!\Selector31~0_combout  & (\Selector27~1_combout  & (\ShiftLeft0~67_combout )))

	.dataa(\Selector31~0_combout ),
	.datab(\Selector27~1_combout ),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\Selector26~2_combout ),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~3 .lut_mask = 16'hEAC0;
defparam \Selector26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N10
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// \Selector4~1_combout  = (\Selector0~2_combout  & ((\input_b~18_combout ) # ((\input_a~69_combout )))) # (!\Selector0~2_combout  & (\input_b~18_combout  & (\Selector0~3_combout  & \input_a~69_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(input_b6),
	.datac(\Selector0~3_combout ),
	.datad(input_a4),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'hEA88;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N26
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// \Selector4~2_combout  = (!\input_b~77_combout  & (\Selector0~0_combout  & (!\ShiftLeft0~24_combout  & !\input_b~79_combout )))

	.dataa(input_b31),
	.datab(\Selector0~0_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(input_b33),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'h0004;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N12
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\input_b~85_combout  & ((\input_a~83_combout ))) # (!\input_b~85_combout  & (\input_a~81_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a10),
	.datad(input_a11),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N26
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\input_b~85_combout  & (\input_a~79_combout )) # (!\input_b~85_combout  & ((\input_a~77_combout )))

	.dataa(input_a9),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a8),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N16
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\input_b~83_combout  & (\ShiftLeft0~64_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~56_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftLeft0~64_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N28
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\input_b~85_combout  & (\input_a~107_combout )) # (!\input_b~85_combout  & ((\input_a~104_combout )))

	.dataa(input_a21),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a20),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N20
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\input_b~83_combout  & (\ShiftLeft0~51_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~68_combout )))

	.dataa(\ShiftLeft0~51_combout ),
	.datab(gnd),
	.datac(input_b37),
	.datad(\ShiftLeft0~68_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N28
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & ((\ShiftLeft0~76_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~80_combout ))))

	.dataa(input_b35),
	.datab(\ShiftLeft0~80_combout ),
	.datac(input_b33),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'h0E04;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\ShiftLeft0~81_combout ) # ((!\input_b~81_combout  & (\input_b~79_combout  & \ShiftLeft0~23_combout )))

	.dataa(input_b35),
	.datab(input_b33),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hFF40;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N28
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\input_b~85_combout  & (\input_a~71_combout )) # (!\input_b~85_combout  & ((\input_a~69_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a5),
	.datad(input_a4),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N12
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\input_b~85_combout  & (\input_a~75_combout )) # (!\input_b~85_combout  & ((\input_a~73_combout )))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a7),
	.datad(input_a6),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N30
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\input_b~83_combout  & ((\ShiftLeft0~57_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~55_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~55_combout ),
	.datac(input_b37),
	.datad(\ShiftLeft0~57_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N24
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\input_b~85_combout  & ((\input_a~91_combout ))) # (!\input_b~85_combout  & (\input_a~89_combout ))

	.dataa(input_a14),
	.datab(input_a15),
	.datac(input_b39),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hCACA;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N28
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\input_b~85_combout  & (\input_a~87_combout )) # (!\input_b~85_combout  & ((\input_a~85_combout )))

	.dataa(input_a13),
	.datab(gnd),
	.datac(input_b39),
	.datad(input_a12),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N30
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\input_b~83_combout  & (\ShiftLeft0~61_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~63_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~61_combout ),
	.datac(input_b37),
	.datad(\ShiftLeft0~63_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N14
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\input_b~85_combout  & ((\input_a~101_combout ))) # (!\input_b~85_combout  & (\input_a~98_combout ))

	.dataa(input_b39),
	.datab(gnd),
	.datac(input_a18),
	.datad(input_a19),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N18
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\input_b~85_combout  & ((\input_a~95_combout ))) # (!\input_b~85_combout  & (\input_a~93_combout ))

	.dataa(gnd),
	.datab(input_a16),
	.datac(input_b39),
	.datad(input_a17),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N0
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\input_b~83_combout  & (\ShiftLeft0~69_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~60_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~69_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N8
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\input_b~81_combout  & ((\ShiftLeft0~83_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~84_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftLeft0~84_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N12
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// \Selector4~3_combout  = (\Selector7~5_combout  & (!\Selector7~13_combout )) # (!\Selector7~5_combout  & ((\Selector7~13_combout  & ((\ShiftLeft0~85_combout ))) # (!\Selector7~13_combout  & (\ShiftLeft0~86_combout ))))

	.dataa(\Selector7~5_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\ShiftLeft0~86_combout ),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'h7632;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N10
cycloneive_lcell_comb \Selector4~4 (
// Equation(s):
// \Selector4~4_combout  = (\Selector7~5_combout  & ((\Selector4~3_combout  & (\ShiftLeft0~79_combout )) # (!\Selector4~3_combout  & ((\ShiftLeft0~82_combout ))))) # (!\Selector7~5_combout  & (((\Selector4~3_combout ))))

	.dataa(\Selector7~5_combout ),
	.datab(\ShiftLeft0~79_combout ),
	.datac(\ShiftLeft0~82_combout ),
	.datad(\Selector4~3_combout ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~4 .lut_mask = 16'hDDA0;
defparam \Selector4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N4
cycloneive_lcell_comb \Selector4~5 (
// Equation(s):
// \Selector4~5_combout  = (\Selector7~4_combout  & ((\Selector4~4_combout ) # ((\ShiftRight0~30_combout  & \Selector4~2_combout )))) # (!\Selector7~4_combout  & (\ShiftRight0~30_combout  & (\Selector4~2_combout )))

	.dataa(\Selector7~4_combout ),
	.datab(\ShiftRight0~30_combout ),
	.datac(\Selector4~2_combout ),
	.datad(\Selector4~4_combout ),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~5 .lut_mask = 16'hEAC0;
defparam \Selector4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N26
cycloneive_lcell_comb \Selector4~6 (
// Equation(s):
// \Selector4~6_combout  = (\Selector4~1_combout ) # ((\Selector4~5_combout ) # ((\Selector0~7_combout  & \Add1~54_combout )))

	.dataa(\Selector4~1_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector4~5_combout ),
	.datad(\Add1~54_combout ),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~6 .lut_mask = 16'hFEFA;
defparam \Selector4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N0
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// \Selector4~0_combout  = (\input_a~69_combout  & (!\input_b~18_combout  & (\Selector0~4_combout ))) # (!\input_a~69_combout  & ((\input_b~18_combout  & (\Selector0~4_combout )) # (!\input_b~18_combout  & ((\Selector0~5_combout )))))

	.dataa(input_a4),
	.datab(input_b6),
	.datac(\Selector0~4_combout ),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'h7160;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N30
cycloneive_lcell_comb \Selector16~9 (
// Equation(s):
// \Selector16~9_combout  = (\Selector0~14_combout  & (!\input_b~77_combout  & (!\ShiftLeft0~20_combout  & !\ShiftLeft0~16_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(input_b31),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~9 .lut_mask = 16'h0002;
defparam \Selector16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N12
cycloneive_lcell_comb \Selector8~2 (
// Equation(s):
// \Selector8~2_combout  = (\input_b~81_combout  & (\ShiftLeft0~80_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~83_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~80_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~2 .lut_mask = 16'hF5A0;
defparam \Selector8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (\input_b~79_combout  & (\ShiftLeft0~77_combout )) # (!\input_b~79_combout  & ((\Selector8~2_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~77_combout ),
	.datac(\Selector8~2_combout ),
	.datad(input_b33),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N4
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\input_b~81_combout ) # ((\input_b~85_combout ) # ((\input_b~83_combout ) # (\input_b~79_combout )))

	.dataa(input_b35),
	.datab(input_b39),
	.datac(input_b37),
	.datad(input_b33),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N12
cycloneive_lcell_comb \Selector16~2 (
// Equation(s):
// \Selector16~2_combout  = (\input_b~77_combout  & (ALUOP_ID_0 & \Selector15~0_combout ))

	.dataa(gnd),
	.datab(input_b31),
	.datac(ALUOP_ID_0),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~2 .lut_mask = 16'hC000;
defparam \Selector16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N4
cycloneive_lcell_comb \Selector16~1 (
// Equation(s):
// \Selector16~1_combout  = (\Selector15~3_combout  & ((\input_b~81_combout  & (\ShiftRight0~29_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~31_combout )))))

	.dataa(\ShiftRight0~29_combout ),
	.datab(input_b35),
	.datac(\ShiftRight0~31_combout ),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~1 .lut_mask = 16'hB800;
defparam \Selector16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N22
cycloneive_lcell_comb \Selector16~3 (
// Equation(s):
// \Selector16~3_combout  = (\Selector16~1_combout ) # ((!\ShiftLeft0~87_combout  & (\Selector16~2_combout  & \input_a~61_combout )))

	.dataa(\ShiftLeft0~87_combout ),
	.datab(\Selector16~2_combout ),
	.datac(input_a),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~3 .lut_mask = 16'hFF40;
defparam \Selector16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N26
cycloneive_lcell_comb \Selector16~4 (
// Equation(s):
// \Selector16~4_combout  = (\input_a~93_combout  & (((!\input_b~54_combout  & \Selector0~10_combout )))) # (!\input_a~93_combout  & ((\input_b~54_combout  & ((\Selector0~10_combout ))) # (!\input_b~54_combout  & (\Selector0~11_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(input_a16),
	.datac(input_b18),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~4 .lut_mask = 16'h3E02;
defparam \Selector16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N2
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\input_b~83_combout  & (\ShiftRight0~25_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~7_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~25_combout ),
	.datad(\ShiftRight0~7_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N30
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\input_b~81_combout  & ((\ShiftRight0~32_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~35_combout ))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftRight0~35_combout ),
	.datad(\ShiftRight0~32_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hFA50;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N24
cycloneive_lcell_comb \Selector16~5 (
// Equation(s):
// \Selector16~5_combout  = (\Selector0~13_combout  & ((\Add1~30_combout ) # ((\Selector0~12_combout  & \Add0~30_combout )))) # (!\Selector0~13_combout  & (((\Selector0~12_combout  & \Add0~30_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Add1~30_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add0~30_combout ),
	.cin(gnd),
	.combout(\Selector16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~5 .lut_mask = 16'hF888;
defparam \Selector16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N22
cycloneive_lcell_comb \Selector16~7 (
// Equation(s):
// \Selector16~7_combout  = (\Selector16~6_combout ) # ((\Selector16~5_combout ) # ((\Selector0~8_combout  & \input_b~54_combout )))

	.dataa(\Selector16~6_combout ),
	.datab(\Selector0~8_combout ),
	.datac(input_b18),
	.datad(\Selector16~5_combout ),
	.cin(gnd),
	.combout(\Selector16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~7 .lut_mask = 16'hFFEA;
defparam \Selector16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N28
cycloneive_lcell_comb \Selector16~8 (
// Equation(s):
// \Selector16~8_combout  = (\Selector16~4_combout ) # ((\Selector16~7_combout ) # ((\Selector16~0_combout  & \ShiftRight0~71_combout )))

	.dataa(\Selector16~4_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\ShiftRight0~71_combout ),
	.datad(\Selector16~7_combout ),
	.cin(gnd),
	.combout(\Selector16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~8 .lut_mask = 16'hFFEA;
defparam \Selector16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N22
cycloneive_lcell_comb \Selector7~8 (
// Equation(s):
// \Selector7~8_combout  = (\Selector0~2_combout  & (((\input_a~75_combout ) # (\input_b~27_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\input_a~75_combout  & \input_b~27_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(input_a7),
	.datad(input_b9),
	.cin(gnd),
	.combout(\Selector7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~8 .lut_mask = 16'hEAA0;
defparam \Selector7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N0
cycloneive_lcell_comb \Selector7~6 (
// Equation(s):
// \Selector7~6_combout  = (\input_a~75_combout  & (\Selector0~4_combout  & ((!\input_b~27_combout )))) # (!\input_a~75_combout  & ((\input_b~27_combout  & (\Selector0~4_combout )) # (!\input_b~27_combout  & ((\Selector0~5_combout )))))

	.dataa(input_a7),
	.datab(\Selector0~4_combout ),
	.datac(\Selector0~5_combout ),
	.datad(input_b9),
	.cin(gnd),
	.combout(\Selector7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~6 .lut_mask = 16'h44D8;
defparam \Selector7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N30
cycloneive_lcell_comb \Selector7~7 (
// Equation(s):
// \Selector7~7_combout  = (Add03 & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add1~48_combout )))) # (!Add03 & (\Selector0~7_combout  & ((\Add1~48_combout ))))

	.dataa(Add03),
	.datab(\Selector0~7_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add1~48_combout ),
	.cin(gnd),
	.combout(\Selector7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~7 .lut_mask = 16'hECA0;
defparam \Selector7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N18
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\input_b~85_combout  & ((\input_a~77_combout ))) # (!\input_b~85_combout  & (\input_a~75_combout ))

	.dataa(input_a7),
	.datab(input_b39),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hE2E2;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N28
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\input_b~85_combout  & ((\input_a~81_combout ))) # (!\input_b~85_combout  & (\input_a~79_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a9),
	.datad(input_a10),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N4
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\input_b~83_combout  & ((\ShiftLeft0~26_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~27_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~27_combout ),
	.datac(input_b37),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N16
cycloneive_lcell_comb \Selector7~9 (
// Equation(s):
// \Selector7~9_combout  = (\Selector7~13_combout  & (\Selector7~5_combout )) # (!\Selector7~13_combout  & ((\Selector7~5_combout  & ((\ShiftLeft0~35_combout ))) # (!\Selector7~5_combout  & (\ShiftLeft0~28_combout ))))

	.dataa(\Selector7~13_combout ),
	.datab(\Selector7~5_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\Selector7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~9 .lut_mask = 16'hDC98;
defparam \Selector7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N30
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\input_b~83_combout  & ((\input_b~85_combout  & ((\input_a~134_combout ))) # (!\input_b~85_combout  & (\input_a~131_combout ))))

	.dataa(input_b37),
	.datab(input_a29),
	.datac(input_a30),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hA088;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N10
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\ShiftLeft0~37_combout ) # ((!\input_b~83_combout  & \ShiftLeft0~38_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N26
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (!\input_b~83_combout  & (\input_b~79_combout  & (!\input_b~81_combout  & !\input_b~85_combout )))

	.dataa(input_b37),
	.datab(input_b33),
	.datac(input_b35),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'h0004;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\input_a~137_combout  & ((\ShiftLeft0~78_combout ) # ((\ShiftLeft0~103_combout  & \ShiftLeft0~43_combout )))) # (!\input_a~137_combout  & (\ShiftLeft0~103_combout  & (\ShiftLeft0~43_combout )))

	.dataa(input_a31),
	.datab(\ShiftLeft0~103_combout ),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~78_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N16
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\ShiftLeft0~90_combout ) # ((\input_b~81_combout  & (!\input_b~79_combout  & \ShiftLeft0~39_combout )))

	.dataa(input_b35),
	.datab(input_b33),
	.datac(\ShiftLeft0~39_combout ),
	.datad(\ShiftLeft0~90_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N18
cycloneive_lcell_comb \Selector7~10 (
// Equation(s):
// \Selector7~10_combout  = (\Selector7~9_combout  & (((\ShiftLeft0~91_combout ) # (!\Selector7~13_combout )))) # (!\Selector7~9_combout  & (\ShiftLeft0~89_combout  & ((\Selector7~13_combout ))))

	.dataa(\ShiftLeft0~89_combout ),
	.datab(\Selector7~9_combout ),
	.datac(\ShiftLeft0~91_combout ),
	.datad(\Selector7~13_combout ),
	.cin(gnd),
	.combout(\Selector7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~10 .lut_mask = 16'hE2CC;
defparam \Selector7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N20
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\input_b~85_combout  & ((\input_a~73_combout ))) # (!\input_b~85_combout  & (\input_a~75_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a7),
	.datad(input_a6),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hFC30;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N30
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\input_b~85_combout  & ((\input_a~69_combout ))) # (!\input_b~85_combout  & (\input_a~71_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_a5),
	.datad(input_a4),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hFC30;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N18
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\input_b~83_combout  & ((\ShiftRight0~54_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~55_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~55_combout ),
	.datac(\ShiftRight0~54_combout ),
	.datad(input_b37),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N14
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\input_b~81_combout  & (\ShiftRight0~40_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~56_combout )))

	.dataa(\ShiftRight0~40_combout ),
	.datab(input_b35),
	.datac(gnd),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hBB88;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N24
cycloneive_lcell_comb \Selector7~11 (
// Equation(s):
// \Selector7~11_combout  = (\Selector7~4_combout  & ((\Selector7~10_combout ) # ((\Selector4~2_combout  & \ShiftRight0~77_combout )))) # (!\Selector7~4_combout  & (((\Selector4~2_combout  & \ShiftRight0~77_combout ))))

	.dataa(\Selector7~4_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\Selector4~2_combout ),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\Selector7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~11 .lut_mask = 16'hF888;
defparam \Selector7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N12
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// \Selector6~0_combout  = (\input_b~24_combout  & (((!\input_a~73_combout  & \Selector0~4_combout )))) # (!\input_b~24_combout  & ((\input_a~73_combout  & ((\Selector0~4_combout ))) # (!\input_a~73_combout  & (\Selector0~5_combout ))))

	.dataa(input_b8),
	.datab(\Selector0~5_combout ),
	.datac(input_a6),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'h5E04;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N14
cycloneive_lcell_comb \Selector6~2 (
// Equation(s):
// \Selector6~2_combout  = (\input_b~24_combout  & ((\Selector0~2_combout ) # ((\Selector0~3_combout  & \input_a~73_combout )))) # (!\input_b~24_combout  & (((\input_a~73_combout  & \Selector0~2_combout ))))

	.dataa(input_b8),
	.datab(\Selector0~3_combout ),
	.datac(input_a6),
	.datad(\Selector0~2_combout ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~2 .lut_mask = 16'hFA80;
defparam \Selector6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N26
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\input_b~83_combout  & (\ShiftLeft0~56_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~57_combout )))

	.dataa(\ShiftLeft0~56_combout ),
	.datab(gnd),
	.datac(input_b37),
	.datad(\ShiftLeft0~57_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N30
cycloneive_lcell_comb \Selector6~3 (
// Equation(s):
// \Selector6~3_combout  = (\Selector7~13_combout  & ((\ShiftLeft0~92_combout ) # ((\Selector7~5_combout )))) # (!\Selector7~13_combout  & (((!\Selector7~5_combout  & \ShiftLeft0~58_combout ))))

	.dataa(\ShiftLeft0~92_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\Selector7~5_combout ),
	.datad(\ShiftLeft0~58_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~3 .lut_mask = 16'hCBC8;
defparam \Selector6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N24
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\input_b~83_combout  & ((\ShiftLeft0~63_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~64_combout ))

	.dataa(\ShiftLeft0~64_combout ),
	.datab(gnd),
	.datac(input_b37),
	.datad(\ShiftLeft0~63_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N20
cycloneive_lcell_comb \Selector6~4 (
// Equation(s):
// \Selector6~4_combout  = (\Selector7~5_combout  & ((\Selector6~3_combout  & (\ShiftLeft0~54_combout )) # (!\Selector6~3_combout  & ((\ShiftLeft0~65_combout ))))) # (!\Selector7~5_combout  & (((\Selector6~3_combout ))))

	.dataa(\ShiftLeft0~54_combout ),
	.datab(\Selector7~5_combout ),
	.datac(\Selector6~3_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~4 .lut_mask = 16'hBCB0;
defparam \Selector6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N10
cycloneive_lcell_comb \Selector6~5 (
// Equation(s):
// \Selector6~5_combout  = (\Selector4~2_combout  & ((\ShiftRight0~20_combout ) # ((\Selector7~4_combout  & \Selector6~4_combout )))) # (!\Selector4~2_combout  & (\Selector7~4_combout  & ((\Selector6~4_combout ))))

	.dataa(\Selector4~2_combout ),
	.datab(\Selector7~4_combout ),
	.datac(\ShiftRight0~20_combout ),
	.datad(\Selector6~4_combout ),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~5 .lut_mask = 16'hECA0;
defparam \Selector6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N12
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// \Selector6~1_combout  = (Add04 & ((\Selector0~6_combout ) # ((\Add1~50_combout  & \Selector0~7_combout )))) # (!Add04 & (((\Add1~50_combout  & \Selector0~7_combout ))))

	.dataa(Add04),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~50_combout ),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'hF888;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N10
cycloneive_lcell_comb \Selector29~2 (
// Equation(s):
// \Selector29~2_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~131_combout ))

	.dataa(gnd),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(input_a29),
	.cin(gnd),
	.combout(\Selector29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~2 .lut_mask = 16'hFCCC;
defparam \Selector29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N16
cycloneive_lcell_comb \Selector29~3 (
// Equation(s):
// \Selector29~3_combout  = (\input_b~81_combout  & ((\Selector29~2_combout ) # ((!\input_a~131_combout  & \Selector0~10_combout )))) # (!\input_b~81_combout  & (\input_a~131_combout  & (\Selector0~10_combout )))

	.dataa(input_b35),
	.datab(input_a29),
	.datac(\Selector0~10_combout ),
	.datad(\Selector29~2_combout ),
	.cin(gnd),
	.combout(\Selector29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~3 .lut_mask = 16'hEA60;
defparam \Selector29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N8
cycloneive_lcell_comb \Selector29~4 (
// Equation(s):
// \Selector29~4_combout  = (\Selector0~12_combout  & ((\Add0~4_combout ) # ((\Selector0~13_combout  & \Add1~4_combout )))) # (!\Selector0~12_combout  & (\Selector0~13_combout  & ((\Add1~4_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add0~4_combout ),
	.datad(\Add1~4_combout ),
	.cin(gnd),
	.combout(\Selector29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~4 .lut_mask = 16'hECA0;
defparam \Selector29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \Selector29~5 (
// Equation(s):
// \Selector29~5_combout  = (\Selector0~11_combout  & (!\input_b~80_combout  & ((!Result_EX_2) # (!\input_b~1_combout ))))

	.dataa(input_b),
	.datab(\Selector0~11_combout ),
	.datac(Result_EX_2),
	.datad(input_b34),
	.cin(gnd),
	.combout(\Selector29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~5 .lut_mask = 16'h004C;
defparam \Selector29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N30
cycloneive_lcell_comb \Selector29~6 (
// Equation(s):
// \Selector29~6_combout  = (\Selector29~4_combout ) # ((\input_a~131_combout  & (\Selector0~8_combout )) # (!\input_a~131_combout  & ((\Selector29~5_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(input_a29),
	.datac(\Selector29~4_combout ),
	.datad(\Selector29~5_combout ),
	.cin(gnd),
	.combout(\Selector29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~6 .lut_mask = 16'hFBF8;
defparam \Selector29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N2
cycloneive_lcell_comb \Selector29~7 (
// Equation(s):
// \Selector29~7_combout  = (\Selector29~3_combout ) # ((\Selector29~6_combout ) # ((\ShiftLeft0~73_combout  & \Selector28~6_combout )))

	.dataa(\Selector29~3_combout ),
	.datab(\Selector29~6_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~7 .lut_mask = 16'hFEEE;
defparam \Selector29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N4
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\input_b~85_combout  & (\input_a~98_combout )) # (!\input_b~85_combout  & ((\input_a~101_combout )))

	.dataa(gnd),
	.datab(input_a18),
	.datac(input_b39),
	.datad(input_a19),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N18
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (\input_b~85_combout  & ((\input_a~104_combout ))) # (!\input_b~85_combout  & (\input_a~107_combout ))

	.dataa(input_a21),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a20),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'hEE22;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N22
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\input_b~83_combout  & (\ShiftRight0~45_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~48_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~45_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N12
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\input_b~81_combout  & (\ShiftRight0~64_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~62_combout )))

	.dataa(\ShiftRight0~64_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~62_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N8
cycloneive_lcell_comb \Selector29~8 (
// Equation(s):
// \Selector29~8_combout  = (\Selector3~1_combout  & (((!\ShiftLeft0~103_combout )))) # (!\Selector3~1_combout  & ((\ShiftLeft0~103_combout  & (\ShiftRight0~80_combout )) # (!\ShiftLeft0~103_combout  & ((\ShiftRight0~66_combout )))))

	.dataa(\ShiftRight0~80_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\ShiftLeft0~103_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\Selector29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~8 .lut_mask = 16'h2F2C;
defparam \Selector29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N2
cycloneive_lcell_comb \Selector29~9 (
// Equation(s):
// \Selector29~9_combout  = (\Selector3~1_combout  & ((\Selector29~8_combout  & ((\ShiftRight0~81_combout ))) # (!\Selector29~8_combout  & (\ShiftRight0~52_combout )))) # (!\Selector3~1_combout  & (((\Selector29~8_combout ))))

	.dataa(\Selector3~1_combout ),
	.datab(\ShiftRight0~52_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(\Selector29~8_combout ),
	.cin(gnd),
	.combout(\Selector29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~9 .lut_mask = 16'hF588;
defparam \Selector29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N22
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\input_b~83_combout  & ((\ShiftRight0~39_combout ))) # (!\input_b~83_combout  & (\ShiftRight0~54_combout ))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftRight0~54_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hFA50;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N6
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\input_b~81_combout  & (!\input_b~83_combout  & ((\ShiftRight0~38_combout )))) # (!\input_b~81_combout  & (((\ShiftRight0~67_combout ))))

	.dataa(input_b37),
	.datab(input_b35),
	.datac(\ShiftRight0~67_combout ),
	.datad(\ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'h7430;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y30_N10
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\input_b~83_combout  & (\ShiftRight0~55_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~57_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~55_combout ),
	.datac(\ShiftRight0~57_combout ),
	.datad(input_b37),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N24
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// \Selector21~0_combout  = (\input_b~81_combout  & (\ShiftRight0~68_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~63_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftRight0~68_combout ),
	.datad(\ShiftRight0~63_combout ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hF5A0;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N6
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\input_b~79_combout  & (\ShiftRight0~78_combout )) # (!\input_b~79_combout  & ((\Selector21~0_combout )))

	.dataa(gnd),
	.datab(input_b33),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N8
cycloneive_lcell_comb \Selector29~1 (
// Equation(s):
// \Selector29~1_combout  = (\input_b~77_combout  & (ALUOP_ID_0 & (\ShiftRight0~79_combout  & \Selector15~0_combout )))

	.dataa(input_b31),
	.datab(ALUOP_ID_0),
	.datac(\ShiftRight0~79_combout ),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~1 .lut_mask = 16'h8000;
defparam \Selector29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N16
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\input_b~81_combout  & ((\ShiftLeft0~46_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~32_combout ))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N12
cycloneive_lcell_comb \Selector15~13 (
// Equation(s):
// \Selector15~13_combout  = (!\ShiftLeft0~24_combout  & (\halt_reg~10_combout  & (!ALUOP_ID_0 & !\Selector15~2_combout )))

	.dataa(\ShiftLeft0~24_combout ),
	.datab(halt_reg),
	.datac(ALUOP_ID_0),
	.datad(\Selector15~2_combout ),
	.cin(gnd),
	.combout(\Selector15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~13 .lut_mask = 16'h0004;
defparam \Selector15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N30
cycloneive_lcell_comb \Selector15~9 (
// Equation(s):
// \Selector15~9_combout  = (\input_b~51_combout  & (\Selector0~10_combout  & (!\input_a~91_combout ))) # (!\input_b~51_combout  & ((\input_a~91_combout  & (\Selector0~10_combout )) # (!\input_a~91_combout  & ((\Selector0~11_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(input_b17),
	.datac(input_a15),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~9 .lut_mask = 16'h2B28;
defparam \Selector15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N18
cycloneive_lcell_comb \Selector15~11 (
// Equation(s):
// \Selector15~11_combout  = (\input_b~51_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~91_combout )))) # (!\input_b~51_combout  & (((\Selector0~8_combout  & \input_a~91_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(input_b17),
	.datac(\Selector0~8_combout ),
	.datad(input_a15),
	.cin(gnd),
	.combout(\Selector15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~11 .lut_mask = 16'hF8C0;
defparam \Selector15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N4
cycloneive_lcell_comb \Selector15~10 (
// Equation(s):
// \Selector15~10_combout  = (\Add1~32_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add0~32_combout )))) # (!\Add1~32_combout  & (\Selector0~12_combout  & (\Add0~32_combout )))

	.dataa(\Add1~32_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~32_combout ),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~10 .lut_mask = 16'hEAC0;
defparam \Selector15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N20
cycloneive_lcell_comb \Selector15~8 (
// Equation(s):
// \Selector15~8_combout  = (\Selector15~1_combout  & ((\input_b~79_combout  & ((\ShiftRight0~77_combout ))) # (!\input_b~79_combout  & (\Selector23~1_combout ))))

	.dataa(\Selector23~1_combout ),
	.datab(\Selector15~1_combout ),
	.datac(input_b33),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\Selector15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~8 .lut_mask = 16'hC808;
defparam \Selector15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N28
cycloneive_lcell_comb \Selector15~12 (
// Equation(s):
// \Selector15~12_combout  = (\Selector15~9_combout ) # ((\Selector15~11_combout ) # ((\Selector15~10_combout ) # (\Selector15~8_combout )))

	.dataa(\Selector15~9_combout ),
	.datab(\Selector15~11_combout ),
	.datac(\Selector15~10_combout ),
	.datad(\Selector15~8_combout ),
	.cin(gnd),
	.combout(\Selector15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~12 .lut_mask = 16'hFFFE;
defparam \Selector15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N26
cycloneive_lcell_comb \Selector15~4 (
// Equation(s):
// \Selector15~4_combout  = (\input_b~79_combout  & (!ALUOP_ID_0 & (!\input_b~77_combout  & \Selector15~0_combout )))

	.dataa(input_b33),
	.datab(ALUOP_ID_0),
	.datac(input_b31),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~4 .lut_mask = 16'h0200;
defparam \Selector15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N8
cycloneive_lcell_comb \Selector15~5 (
// Equation(s):
// \Selector15~5_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & ((\ShiftLeft0~39_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~43_combout ),
	.datab(\Selector15~4_combout ),
	.datac(\ShiftLeft0~39_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\Selector15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~5 .lut_mask = 16'hC088;
defparam \Selector15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N0
cycloneive_lcell_comb \Selector15~6 (
// Equation(s):
// \Selector15~6_combout  = (!ALUOP_ID_0 & (\input_b~77_combout  & \Selector15~0_combout ))

	.dataa(gnd),
	.datab(ALUOP_ID_0),
	.datac(input_b31),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~6 .lut_mask = 16'h3000;
defparam \Selector15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N26
cycloneive_lcell_comb \Selector15~7 (
// Equation(s):
// \Selector15~7_combout  = (\Selector15~5_combout ) # ((\input_a~137_combout  & (!\ShiftLeft0~87_combout  & \Selector15~6_combout )))

	.dataa(input_a31),
	.datab(\ShiftLeft0~87_combout ),
	.datac(\Selector15~5_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~7 .lut_mask = 16'hF2F0;
defparam \Selector15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N6
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (\input_b~21_combout  & (((!\input_a~71_combout  & \Selector0~4_combout )))) # (!\input_b~21_combout  & ((\input_a~71_combout  & ((\Selector0~4_combout ))) # (!\input_a~71_combout  & (\Selector0~5_combout ))))

	.dataa(input_b7),
	.datab(\Selector0~5_combout ),
	.datac(input_a5),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'h5E04;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N2
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// \Selector5~2_combout  = (\Selector0~2_combout  & (((\input_a~71_combout ) # (\input_b~21_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\input_a~71_combout  & \input_b~21_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(input_a5),
	.datad(input_b7),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hEAA0;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N14
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (\input_b~83_combout  & ((\ShiftLeft0~42_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~44_combout ))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N10
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (!\input_b~79_combout  & ((\input_b~81_combout  & (\ShiftLeft0~74_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~98_combout )))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(input_b35),
	.datac(input_b33),
	.datad(\ShiftLeft0~98_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'h0B08;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N8
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (\ShiftLeft0~99_combout ) # ((\ShiftLeft0~73_combout  & (!\input_b~81_combout  & \input_b~79_combout )))

	.dataa(\ShiftLeft0~73_combout ),
	.datab(input_b35),
	.datac(input_b33),
	.datad(\ShiftLeft0~99_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N24
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (\input_b~83_combout  & ((\ShiftLeft0~27_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~25_combout ))

	.dataa(\ShiftLeft0~25_combout ),
	.datab(\ShiftLeft0~27_combout ),
	.datac(input_b37),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hCACA;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N18
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (\input_b~83_combout  & ((\ShiftLeft0~34_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~26_combout ))

	.dataa(input_b37),
	.datab(\ShiftLeft0~26_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N28
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (\Selector7~13_combout  & (((\Selector7~5_combout )))) # (!\Selector7~13_combout  & ((\Selector7~5_combout  & ((\ShiftLeft0~96_combout ))) # (!\Selector7~5_combout  & (\ShiftLeft0~97_combout ))))

	.dataa(\Selector7~13_combout ),
	.datab(\ShiftLeft0~97_combout ),
	.datac(\Selector7~5_combout ),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'hF4A4;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N6
cycloneive_lcell_comb \Selector5~4 (
// Equation(s):
// \Selector5~4_combout  = (\Selector7~13_combout  & ((\Selector5~3_combout  & ((\ShiftLeft0~100_combout ))) # (!\Selector5~3_combout  & (\ShiftLeft0~95_combout )))) # (!\Selector7~13_combout  & (((\Selector5~3_combout ))))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(\Selector7~13_combout ),
	.datac(\ShiftLeft0~100_combout ),
	.datad(\Selector5~3_combout ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~4 .lut_mask = 16'hF388;
defparam \Selector5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N8
cycloneive_lcell_comb \Selector5~5 (
// Equation(s):
// \Selector5~5_combout  = (\Selector7~4_combout  & ((\Selector5~4_combout ) # ((\ShiftRight0~78_combout  & \Selector4~2_combout )))) # (!\Selector7~4_combout  & (\ShiftRight0~78_combout  & (\Selector4~2_combout )))

	.dataa(\Selector7~4_combout ),
	.datab(\ShiftRight0~78_combout ),
	.datac(\Selector4~2_combout ),
	.datad(\Selector5~4_combout ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~5 .lut_mask = 16'hEAC0;
defparam \Selector5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y30_N28
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// \Selector5~1_combout  = (Add05 & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add1~52_combout )))) # (!Add05 & (((\Selector0~7_combout  & \Add1~52_combout ))))

	.dataa(Add05),
	.datab(\Selector0~6_combout ),
	.datac(\Selector0~7_combout ),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'hF888;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((!\input_a~137_combout  & \input_b~85_combout ))

	.dataa(input_a31),
	.datab(input_b39),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\input_a~134_combout  & ((!\LessThan0~1_cout ) # (!\input_b~83_combout ))) # (!\input_a~134_combout  & (!\input_b~83_combout  & !\LessThan0~1_cout )))

	.dataa(input_a30),
	.datab(input_b37),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\input_b~81_combout  & ((!\LessThan0~3_cout ) # (!\input_a~131_combout ))) # (!\input_b~81_combout  & (!\input_a~131_combout  & !\LessThan0~3_cout )))

	.dataa(input_b35),
	.datab(input_a29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\input_a~128_combout  & ((!\LessThan0~5_cout ) # (!\input_b~79_combout ))) # (!\input_a~128_combout  & (!\input_b~79_combout  & !\LessThan0~5_cout )))

	.dataa(input_a28),
	.datab(input_b33),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\input_a~125_combout  & (\input_b~77_combout  & !\LessThan0~7_cout )) # (!\input_a~125_combout  & ((\input_b~77_combout ) # (!\LessThan0~7_cout ))))

	.dataa(input_a27),
	.datab(input_b31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\input_b~75_combout  & (\input_a~122_combout  & !\LessThan0~9_cout )) # (!\input_b~75_combout  & ((\input_a~122_combout ) # (!\LessThan0~9_cout ))))

	.dataa(input_b29),
	.datab(input_a26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\input_b~73_combout  & ((!\LessThan0~11_cout ) # (!\input_a~119_combout ))) # (!\input_b~73_combout  & (!\input_a~119_combout  & !\LessThan0~11_cout )))

	.dataa(input_b28),
	.datab(input_a25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((\input_b~71_combout  & (\input_a~116_combout  & !\LessThan0~13_cout )) # (!\input_b~71_combout  & ((\input_a~116_combout ) # (!\LessThan0~13_cout ))))

	.dataa(input_b27),
	.datab(input_a24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h004D;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\input_a~113_combout  & (\input_b~69_combout  & !\LessThan0~15_cout )) # (!\input_a~113_combout  & ((\input_b~69_combout ) # (!\LessThan0~15_cout ))))

	.dataa(input_a23),
	.datab(input_b25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((\input_a~110_combout  & ((!\LessThan0~17_cout ) # (!\input_b~67_combout ))) # (!\input_a~110_combout  & (!\input_b~67_combout  & !\LessThan0~17_cout )))

	.dataa(input_a22),
	.datab(input_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\input_a~107_combout  & (\input_b~65_combout  & !\LessThan0~19_cout )) # (!\input_a~107_combout  & ((\input_b~65_combout ) # (!\LessThan0~19_cout ))))

	.dataa(input_a21),
	.datab(input_b23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h004D;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\input_b~63_combout  & (\input_a~104_combout  & !\LessThan0~21_cout )) # (!\input_b~63_combout  & ((\input_a~104_combout ) # (!\LessThan0~21_cout ))))

	.dataa(input_b22),
	.datab(input_a20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((\input_a~101_combout  & (\input_b~61_combout  & !\LessThan0~23_cout )) # (!\input_a~101_combout  & ((\input_b~61_combout ) # (!\LessThan0~23_cout ))))

	.dataa(input_a19),
	.datab(input_b21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\input_a~98_combout  & ((!\LessThan0~25_cout ) # (!\input_b~59_combout ))) # (!\input_a~98_combout  & (!\input_b~59_combout  & !\LessThan0~25_cout )))

	.dataa(input_a18),
	.datab(input_b20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h002B;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\input_b~57_combout  & ((!\LessThan0~27_cout ) # (!\input_a~95_combout ))) # (!\input_b~57_combout  & (!\input_a~95_combout  & !\LessThan0~27_cout )))

	.dataa(input_b19),
	.datab(input_a17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h002B;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\input_b~54_combout  & (\input_a~93_combout  & !\LessThan0~29_cout )) # (!\input_b~54_combout  & ((\input_a~93_combout ) # (!\LessThan0~29_cout ))))

	.dataa(input_b18),
	.datab(input_a16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h004D;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\input_a~91_combout  & (\input_b~51_combout  & !\LessThan0~31_cout )) # (!\input_a~91_combout  & ((\input_b~51_combout ) # (!\LessThan0~31_cout ))))

	.dataa(input_a15),
	.datab(input_b17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\input_a~89_combout  & ((!\LessThan0~33_cout ) # (!\input_b~48_combout ))) # (!\input_a~89_combout  & (!\input_b~48_combout  & !\LessThan0~33_cout )))

	.dataa(input_a14),
	.datab(input_b16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h002B;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\input_b~45_combout  & ((!\LessThan0~35_cout ) # (!\input_a~87_combout ))) # (!\input_b~45_combout  & (!\input_a~87_combout  & !\LessThan0~35_cout )))

	.dataa(input_b15),
	.datab(input_a13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h002B;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((\input_b~42_combout  & (\input_a~85_combout  & !\LessThan0~37_cout )) # (!\input_b~42_combout  & ((\input_a~85_combout ) # (!\LessThan0~37_cout ))))

	.dataa(input_b14),
	.datab(input_a12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h004D;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\input_b~39_combout  & ((!\LessThan0~39_cout ) # (!\input_a~83_combout ))) # (!\input_b~39_combout  & (!\input_a~83_combout  & !\LessThan0~39_cout )))

	.dataa(input_b13),
	.datab(input_a11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h002B;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\input_b~36_combout  & (\input_a~81_combout  & !\LessThan0~41_cout )) # (!\input_b~36_combout  & ((\input_a~81_combout ) # (!\LessThan0~41_cout ))))

	.dataa(input_b12),
	.datab(input_a10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\input_b~33_combout  & ((!\LessThan0~43_cout ) # (!\input_a~79_combout ))) # (!\input_b~33_combout  & (!\input_a~79_combout  & !\LessThan0~43_cout )))

	.dataa(input_b11),
	.datab(input_a9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h002B;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\input_b~30_combout  & (\input_a~77_combout  & !\LessThan0~45_cout )) # (!\input_b~30_combout  & ((\input_a~77_combout ) # (!\LessThan0~45_cout ))))

	.dataa(input_b10),
	.datab(input_a8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h004D;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\input_b~27_combout  & ((!\LessThan0~47_cout ) # (!\input_a~75_combout ))) # (!\input_b~27_combout  & (!\input_a~75_combout  & !\LessThan0~47_cout )))

	.dataa(input_b9),
	.datab(input_a7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\input_a~73_combout  & ((!\LessThan0~49_cout ) # (!\input_b~24_combout ))) # (!\input_a~73_combout  & (!\input_b~24_combout  & !\LessThan0~49_cout )))

	.dataa(input_a6),
	.datab(input_b8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h002B;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\input_b~21_combout  & ((!\LessThan0~51_cout ) # (!\input_a~71_combout ))) # (!\input_b~21_combout  & (!\input_a~71_combout  & !\LessThan0~51_cout )))

	.dataa(input_b7),
	.datab(input_a5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h002B;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\input_b~18_combout  & (\input_a~69_combout  & !\LessThan0~53_cout )) # (!\input_b~18_combout  & ((\input_a~69_combout ) # (!\LessThan0~53_cout ))))

	.dataa(input_b6),
	.datab(input_a4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h004D;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\input_a~67_combout  & (\input_b~15_combout  & !\LessThan0~55_cout )) # (!\input_a~67_combout  & ((\input_b~15_combout ) # (!\LessThan0~55_cout ))))

	.dataa(input_a3),
	.datab(input_b5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\input_b~12_combout  & (\input_a~65_combout  & !\LessThan0~57_cout )) # (!\input_b~12_combout  & ((\input_a~65_combout ) # (!\LessThan0~57_cout ))))

	.dataa(input_b4),
	.datab(input_a2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h004D;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((\input_a~63_combout  & (\input_b~9_combout  & !\LessThan0~59_cout )) # (!\input_a~63_combout  & ((\input_b~9_combout ) # (!\LessThan0~59_cout ))))

	.dataa(input_a1),
	.datab(input_b3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\input_b~6_combout  & (\LessThan0~61_cout  & \input_a~61_combout )) # (!\input_b~6_combout  & ((\LessThan0~61_cout ) # (\input_a~61_combout )))

	.dataa(input_b2),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF550;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N26
cycloneive_lcell_comb \Selector0~16 (
// Equation(s):
// \Selector0~16_combout  = (!ALUOP_ID_2 & (!ALUOP_ID_0 & (ALUOP_ID_1 & ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~16 .lut_mask = 16'h1000;
defparam \Selector0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N6
cycloneive_lcell_comb \Selector31~1 (
// Equation(s):
// \Selector31~1_combout  = (\Selector0~5_combout  & (!\input_a~137_combout  & !\input_b~85_combout ))

	.dataa(gnd),
	.datab(\Selector0~5_combout ),
	.datac(input_a31),
	.datad(input_b39),
	.cin(gnd),
	.combout(\Selector31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~1 .lut_mask = 16'h000C;
defparam \Selector31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N22
cycloneive_lcell_comb \Selector31~9 (
// Equation(s):
// \Selector31~9_combout  = (\Selector0~2_combout  & ((\input_b~84_combout ) # ((\input_b~1_combout  & Result_EX_0))))

	.dataa(\Selector0~2_combout ),
	.datab(input_b38),
	.datac(input_b),
	.datad(Result_EX_0),
	.cin(gnd),
	.combout(\Selector31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~9 .lut_mask = 16'hA888;
defparam \Selector31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((!\input_a~137_combout  & \input_b~85_combout ))

	.dataa(input_a31),
	.datab(input_b39),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0044;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\input_b~83_combout  & (\input_a~134_combout  & !\LessThan1~1_cout )) # (!\input_b~83_combout  & ((\input_a~134_combout ) # (!\LessThan1~1_cout ))))

	.dataa(input_b37),
	.datab(input_a30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h004D;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\input_b~81_combout  & ((!\LessThan1~3_cout ) # (!\input_a~131_combout ))) # (!\input_b~81_combout  & (!\input_a~131_combout  & !\LessThan1~3_cout )))

	.dataa(input_b35),
	.datab(input_a29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h002B;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\input_a~128_combout  & ((!\LessThan1~5_cout ) # (!\input_b~79_combout ))) # (!\input_a~128_combout  & (!\input_b~79_combout  & !\LessThan1~5_cout )))

	.dataa(input_a28),
	.datab(input_b33),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\input_a~125_combout  & (\input_b~77_combout  & !\LessThan1~7_cout )) # (!\input_a~125_combout  & ((\input_b~77_combout ) # (!\LessThan1~7_cout ))))

	.dataa(input_a27),
	.datab(input_b31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\input_a~122_combout  & ((!\LessThan1~9_cout ) # (!\input_b~75_combout ))) # (!\input_a~122_combout  & (!\input_b~75_combout  & !\LessThan1~9_cout )))

	.dataa(input_a26),
	.datab(input_b29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h002B;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\input_a~119_combout  & (\input_b~73_combout  & !\LessThan1~11_cout )) # (!\input_a~119_combout  & ((\input_b~73_combout ) # (!\LessThan1~11_cout ))))

	.dataa(input_a25),
	.datab(input_b28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\input_b~71_combout  & (\input_a~116_combout  & !\LessThan1~13_cout )) # (!\input_b~71_combout  & ((\input_a~116_combout ) # (!\LessThan1~13_cout ))))

	.dataa(input_b27),
	.datab(input_a24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h004D;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\input_a~113_combout  & (\input_b~69_combout  & !\LessThan1~15_cout )) # (!\input_a~113_combout  & ((\input_b~69_combout ) # (!\LessThan1~15_cout ))))

	.dataa(input_a23),
	.datab(input_b25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\input_a~110_combout  & ((!\LessThan1~17_cout ) # (!\input_b~67_combout ))) # (!\input_a~110_combout  & (!\input_b~67_combout  & !\LessThan1~17_cout )))

	.dataa(input_a22),
	.datab(input_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\input_b~65_combout  & ((!\LessThan1~19_cout ) # (!\input_a~107_combout ))) # (!\input_b~65_combout  & (!\input_a~107_combout  & !\LessThan1~19_cout )))

	.dataa(input_b23),
	.datab(input_a21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\input_a~104_combout  & ((!\LessThan1~21_cout ) # (!\input_b~63_combout ))) # (!\input_a~104_combout  & (!\input_b~63_combout  & !\LessThan1~21_cout )))

	.dataa(input_a20),
	.datab(input_b22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h002B;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\input_b~61_combout  & ((!\LessThan1~23_cout ) # (!\input_a~101_combout ))) # (!\input_b~61_combout  & (!\input_a~101_combout  & !\LessThan1~23_cout )))

	.dataa(input_b21),
	.datab(input_a19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h002B;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\input_b~59_combout  & (\input_a~98_combout  & !\LessThan1~25_cout )) # (!\input_b~59_combout  & ((\input_a~98_combout ) # (!\LessThan1~25_cout ))))

	.dataa(input_b20),
	.datab(input_a18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h004D;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\input_b~57_combout  & ((!\LessThan1~27_cout ) # (!\input_a~95_combout ))) # (!\input_b~57_combout  & (!\input_a~95_combout  & !\LessThan1~27_cout )))

	.dataa(input_b19),
	.datab(input_a17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h002B;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((\input_a~93_combout  & ((!\LessThan1~29_cout ) # (!\input_b~54_combout ))) # (!\input_a~93_combout  & (!\input_b~54_combout  & !\LessThan1~29_cout )))

	.dataa(input_a16),
	.datab(input_b18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\input_b~51_combout  & ((!\LessThan1~31_cout ) # (!\input_a~91_combout ))) # (!\input_b~51_combout  & (!\input_a~91_combout  & !\LessThan1~31_cout )))

	.dataa(input_b17),
	.datab(input_a15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\input_a~89_combout  & ((!\LessThan1~33_cout ) # (!\input_b~48_combout ))) # (!\input_a~89_combout  & (!\input_b~48_combout  & !\LessThan1~33_cout )))

	.dataa(input_a14),
	.datab(input_b16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h002B;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\input_b~45_combout  & ((!\LessThan1~35_cout ) # (!\input_a~87_combout ))) # (!\input_b~45_combout  & (!\input_a~87_combout  & !\LessThan1~35_cout )))

	.dataa(input_b15),
	.datab(input_a13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\input_a~85_combout  & ((!\LessThan1~37_cout ) # (!\input_b~42_combout ))) # (!\input_a~85_combout  & (!\input_b~42_combout  & !\LessThan1~37_cout )))

	.dataa(input_a12),
	.datab(input_b14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h002B;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\input_a~83_combout  & (\input_b~39_combout  & !\LessThan1~39_cout )) # (!\input_a~83_combout  & ((\input_b~39_combout ) # (!\LessThan1~39_cout ))))

	.dataa(input_a11),
	.datab(input_b13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\input_b~36_combout  & (\input_a~81_combout  & !\LessThan1~41_cout )) # (!\input_b~36_combout  & ((\input_a~81_combout ) # (!\LessThan1~41_cout ))))

	.dataa(input_b12),
	.datab(input_a10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h004D;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\input_a~79_combout  & (\input_b~33_combout  & !\LessThan1~43_cout )) # (!\input_a~79_combout  & ((\input_b~33_combout ) # (!\LessThan1~43_cout ))))

	.dataa(input_a9),
	.datab(input_b11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h004D;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\input_a~77_combout  & ((!\LessThan1~45_cout ) # (!\input_b~30_combout ))) # (!\input_a~77_combout  & (!\input_b~30_combout  & !\LessThan1~45_cout )))

	.dataa(input_a8),
	.datab(input_b10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h002B;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\input_a~75_combout  & (\input_b~27_combout  & !\LessThan1~47_cout )) # (!\input_a~75_combout  & ((\input_b~27_combout ) # (!\LessThan1~47_cout ))))

	.dataa(input_a7),
	.datab(input_b9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h004D;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\input_b~24_combout  & (\input_a~73_combout  & !\LessThan1~49_cout )) # (!\input_b~24_combout  & ((\input_a~73_combout ) # (!\LessThan1~49_cout ))))

	.dataa(input_b8),
	.datab(input_a6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h004D;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((\input_b~21_combout  & ((!\LessThan1~51_cout ) # (!\input_a~71_combout ))) # (!\input_b~21_combout  & (!\input_a~71_combout  & !\LessThan1~51_cout )))

	.dataa(input_b7),
	.datab(input_a5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h002B;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\input_a~69_combout  & ((!\LessThan1~53_cout ) # (!\input_b~18_combout ))) # (!\input_a~69_combout  & (!\input_b~18_combout  & !\LessThan1~53_cout )))

	.dataa(input_a4),
	.datab(input_b6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h002B;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\input_a~67_combout  & (\input_b~15_combout  & !\LessThan1~55_cout )) # (!\input_a~67_combout  & ((\input_b~15_combout ) # (!\LessThan1~55_cout ))))

	.dataa(input_a3),
	.datab(input_b5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h004D;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\input_b~12_combout  & (\input_a~65_combout  & !\LessThan1~57_cout )) # (!\input_b~12_combout  & ((\input_a~65_combout ) # (!\LessThan1~57_cout ))))

	.dataa(input_b4),
	.datab(input_a2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h004D;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\input_a~63_combout  & (\input_b~9_combout  & !\LessThan1~59_cout )) # (!\input_a~63_combout  & ((\input_b~9_combout ) # (!\LessThan1~59_cout ))))

	.dataa(input_a1),
	.datab(input_b3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\input_a~61_combout  & (\LessThan1~61_cout  & \input_b~6_combout )) # (!\input_a~61_combout  & ((\LessThan1~61_cout ) # (\input_b~6_combout )))

	.dataa(gnd),
	.datab(input_a),
	.datac(gnd),
	.datad(input_b2),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF330;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N28
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (!\input_b~83_combout  & ((\input_b~85_combout  & (\input_a~134_combout )) # (!\input_b~85_combout  & ((\input_a~137_combout )))))

	.dataa(input_b37),
	.datab(input_a30),
	.datac(input_a31),
	.datad(input_b39),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'h4450;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N24
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (!\input_b~81_combout  & ((\ShiftRight0~82_combout ) # ((\ShiftRight0~80_combout  & \input_b~83_combout ))))

	.dataa(\ShiftRight0~80_combout ),
	.datab(\ShiftRight0~82_combout ),
	.datac(input_b37),
	.datad(input_b35),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'h00EC;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N26
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (!\input_b~79_combout  & ((\ShiftRight0~83_combout ) # ((\input_b~81_combout  & \ShiftRight0~53_combout ))))

	.dataa(input_b35),
	.datab(input_b33),
	.datac(\ShiftRight0~53_combout ),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'h3320;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N20
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (!\input_b~77_combout  & ((\ShiftRight0~84_combout ) # ((\ShiftRight0~85_combout  & \input_b~79_combout ))))

	.dataa(\ShiftRight0~85_combout ),
	.datab(input_b31),
	.datac(input_b33),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'h3320;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N8
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (!ALUOP_ID_3 & (!ALUOP_ID_1 & (!ALUOP_ID_0 & !ALUOP_ID_2)))

	.dataa(ALUOP_ID_3),
	.datab(ALUOP_ID_1),
	.datac(ALUOP_ID_0),
	.datad(ALUOP_ID_2),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'h0001;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N8
cycloneive_lcell_comb \Selector31~4 (
// Equation(s):
// \Selector31~4_combout  = (!\ShiftLeft0~87_combout  & (\Selector0~1_combout  & (!\ShiftLeft0~24_combout  & !\input_b~77_combout )))

	.dataa(\ShiftLeft0~87_combout ),
	.datab(\Selector0~1_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(input_b31),
	.cin(gnd),
	.combout(\Selector31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~4 .lut_mask = 16'h0004;
defparam \Selector31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N2
cycloneive_lcell_comb \Selector31~5 (
// Equation(s):
// \Selector31~5_combout  = (\Selector31~4_combout ) # ((\Selector0~2_combout ) # ((\Selector0~3_combout  & \input_b~85_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(input_b39),
	.datac(\Selector31~4_combout ),
	.datad(\Selector0~2_combout ),
	.cin(gnd),
	.combout(\Selector31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~5 .lut_mask = 16'hFFF8;
defparam \Selector31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N20
cycloneive_lcell_comb \Selector31~7 (
// Equation(s):
// \Selector31~7_combout  = (\Selector31~6_combout  & ((\Selector31~0_combout ) # ((\input_a~137_combout  & \Selector31~5_combout )))) # (!\Selector31~6_combout  & (((\input_a~137_combout  & \Selector31~5_combout ))))

	.dataa(\Selector31~6_combout ),
	.datab(\Selector31~0_combout ),
	.datac(input_a31),
	.datad(\Selector31~5_combout ),
	.cin(gnd),
	.combout(\Selector31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~7 .lut_mask = 16'hF888;
defparam \Selector31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N22
cycloneive_lcell_comb \Selector31~8 (
// Equation(s):
// \Selector31~8_combout  = (\Selector31~3_combout ) # ((\Selector31~7_combout ) # ((\Selector31~0_combout  & \ShiftRight0~86_combout )))

	.dataa(\Selector31~3_combout ),
	.datab(\Selector31~0_combout ),
	.datac(\ShiftRight0~86_combout ),
	.datad(\Selector31~7_combout ),
	.cin(gnd),
	.combout(\Selector31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~8 .lut_mask = 16'hFFEA;
defparam \Selector31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N4
cycloneive_lcell_comb \Selector0~17 (
// Equation(s):
// \Selector0~17_combout  = (!ALUOP_ID_2 & (ALUOP_ID_0 & (ALUOP_ID_1 & ALUOP_ID_3)))

	.dataa(ALUOP_ID_2),
	.datab(ALUOP_ID_0),
	.datac(ALUOP_ID_1),
	.datad(ALUOP_ID_3),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~17 .lut_mask = 16'h4000;
defparam \Selector0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N24
cycloneive_lcell_comb \Selector31~10 (
// Equation(s):
// \Selector31~10_combout  = (\Selector31~9_combout ) # ((\Selector31~8_combout ) # ((\LessThan1~62_combout  & \Selector0~17_combout )))

	.dataa(\Selector31~9_combout ),
	.datab(\LessThan1~62_combout ),
	.datac(\Selector31~8_combout ),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~10 .lut_mask = 16'hFEFA;
defparam \Selector31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N22
cycloneive_lcell_comb \Selector11~4 (
// Equation(s):
// \Selector11~4_combout  = (!\input_b~79_combout  & (\input_b~77_combout  & (!ALUOP_ID_0 & \Selector15~0_combout )))

	.dataa(input_b33),
	.datab(input_b31),
	.datac(ALUOP_ID_0),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~4 .lut_mask = 16'h0400;
defparam \Selector11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N30
cycloneive_lcell_comb \Selector11~3 (
// Equation(s):
// \Selector11~3_combout  = (\Add1~40_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add0~40_combout )))) # (!\Add1~40_combout  & (\Selector0~12_combout  & (\Add0~40_combout )))

	.dataa(\Add1~40_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~40_combout ),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~3 .lut_mask = 16'hEAC0;
defparam \Selector11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N10
cycloneive_lcell_comb \Selector11~5 (
// Equation(s):
// \Selector11~5_combout  = (\input_a~83_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_b~39_combout )))) # (!\input_a~83_combout  & (((\Selector0~8_combout  & \input_b~39_combout ))))

	.dataa(input_a11),
	.datab(\Selector0~9_combout ),
	.datac(\Selector0~8_combout ),
	.datad(input_b13),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~5 .lut_mask = 16'hF8A0;
defparam \Selector11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N0
cycloneive_lcell_comb \Selector11~6 (
// Equation(s):
// \Selector11~6_combout  = (\input_a~83_combout  & (\Selector0~10_combout  & ((!\input_b~39_combout )))) # (!\input_a~83_combout  & ((\input_b~39_combout  & (\Selector0~10_combout )) # (!\input_b~39_combout  & ((\Selector0~11_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~11_combout ),
	.datac(input_a11),
	.datad(input_b13),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~6 .lut_mask = 16'h0AAC;
defparam \Selector11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N20
cycloneive_lcell_comb \Selector11~10 (
// Equation(s):
// \Selector11~10_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & (\ShiftLeft0~43_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~46_combout )))))

	.dataa(\ShiftLeft0~43_combout ),
	.datab(input_b35),
	.datac(\Selector15~4_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\Selector11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~10 .lut_mask = 16'hB080;
defparam \Selector11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N0
cycloneive_lcell_comb \Selector11~7 (
// Equation(s):
// \Selector11~7_combout  = (\Selector11~6_combout ) # ((\Selector11~10_combout ) # ((\Selector15~1_combout  & \ShiftRight0~61_combout )))

	.dataa(\Selector15~1_combout ),
	.datab(\Selector11~6_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\Selector11~10_combout ),
	.cin(gnd),
	.combout(\Selector11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~7 .lut_mask = 16'hFFEC;
defparam \Selector11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N28
cycloneive_lcell_comb \Selector11~8 (
// Equation(s):
// \Selector11~8_combout  = (\Selector11~5_combout ) # ((\Selector11~7_combout ) # ((\ShiftLeft0~36_combout  & \Selector15~13_combout )))

	.dataa(\Selector11~5_combout ),
	.datab(\ShiftLeft0~36_combout ),
	.datac(\Selector15~13_combout ),
	.datad(\Selector11~7_combout ),
	.cin(gnd),
	.combout(\Selector11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~8 .lut_mask = 16'hFFEA;
defparam \Selector11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N16
cycloneive_lcell_comb \Selector10~3 (
// Equation(s):
// \Selector10~3_combout  = (\Add1~42_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & Add0)))) # (!\Add1~42_combout  & (((\Selector0~12_combout  & Add0))))

	.dataa(\Add1~42_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(Add0),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~3 .lut_mask = 16'hF888;
defparam \Selector10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y27_N6
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\input_b~83_combout  & (\ShiftLeft0~60_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~61_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~60_combout ),
	.datac(input_b37),
	.datad(\ShiftLeft0~61_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N2
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\input_b~81_combout  & (\ShiftLeft0~62_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~65_combout )))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftLeft0~62_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \Selector10~4 (
// Equation(s):
// \Selector10~4_combout  = (\Selector0~8_combout  & (((\input_a~81_combout ) # (\input_b~36_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\input_a~81_combout  & \input_b~36_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(input_a10),
	.datad(input_b12),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~4 .lut_mask = 16'hECC0;
defparam \Selector10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N6
cycloneive_lcell_comb \Selector10~5 (
// Equation(s):
// \Selector10~5_combout  = (\input_b~36_combout  & (((\Selector0~10_combout  & !\input_a~81_combout )))) # (!\input_b~36_combout  & ((\input_a~81_combout  & ((\Selector0~10_combout ))) # (!\input_a~81_combout  & (\Selector0~11_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(input_b12),
	.datac(\Selector0~10_combout ),
	.datad(input_a10),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~5 .lut_mask = 16'h30E2;
defparam \Selector10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N28
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\input_b~83_combout  & ((\ShiftLeft0~68_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~69_combout ))

	.dataa(\ShiftLeft0~69_combout ),
	.datab(gnd),
	.datac(input_b37),
	.datad(\ShiftLeft0~68_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N6
cycloneive_lcell_comb \Selector10~9 (
// Equation(s):
// \Selector10~9_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & (\ShiftLeft0~52_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~70_combout )))))

	.dataa(\ShiftLeft0~52_combout ),
	.datab(input_b35),
	.datac(\Selector15~4_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\Selector10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~9 .lut_mask = 16'hB080;
defparam \Selector10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N18
cycloneive_lcell_comb \Selector10~6 (
// Equation(s):
// \Selector10~6_combout  = (\Selector10~5_combout ) # ((\Selector10~9_combout ) # ((\Selector15~1_combout  & \ShiftRight0~76_combout )))

	.dataa(\Selector15~1_combout ),
	.datab(\Selector10~5_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\Selector10~9_combout ),
	.cin(gnd),
	.combout(\Selector10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~6 .lut_mask = 16'hFFEC;
defparam \Selector10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N0
cycloneive_lcell_comb \Selector10~7 (
// Equation(s):
// \Selector10~7_combout  = (\Selector10~4_combout ) # ((\Selector10~6_combout ) # ((\Selector15~13_combout  & \ShiftLeft0~66_combout )))

	.dataa(\Selector15~13_combout ),
	.datab(\ShiftLeft0~66_combout ),
	.datac(\Selector10~4_combout ),
	.datad(\Selector10~6_combout ),
	.cin(gnd),
	.combout(\Selector10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~7 .lut_mask = 16'hFFF8;
defparam \Selector10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y27_N10
cycloneive_lcell_comb \Selector21~1 (
// Equation(s):
// \Selector21~1_combout  = (\Selector16~9_combout  & \ShiftLeft0~100_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector16~9_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~1 .lut_mask = 16'hF000;
defparam \Selector21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N28
cycloneive_lcell_comb \Selector21~2 (
// Equation(s):
// \Selector21~2_combout  = (\input_b~65_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~107_combout ))))

	.dataa(input_b23),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(input_a21),
	.cin(gnd),
	.combout(\Selector21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~2 .lut_mask = 16'hA888;
defparam \Selector21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y28_N18
cycloneive_lcell_comb \Selector21~3 (
// Equation(s):
// \Selector21~3_combout  = (\Selector21~2_combout ) # ((\Selector0~10_combout  & (\input_b~65_combout  $ (\input_a~107_combout ))))

	.dataa(input_b23),
	.datab(input_a21),
	.datac(\Selector0~10_combout ),
	.datad(\Selector21~2_combout ),
	.cin(gnd),
	.combout(\Selector21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~3 .lut_mask = 16'hFF60;
defparam \Selector21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N2
cycloneive_lcell_comb \Selector21~7 (
// Equation(s):
// \Selector21~7_combout  = (\Selector21~6_combout ) # ((\Selector21~3_combout ) # ((\Selector16~0_combout  & \ShiftRight0~81_combout )))

	.dataa(\Selector21~6_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector21~3_combout ),
	.datad(\ShiftRight0~81_combout ),
	.cin(gnd),
	.combout(\Selector21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~7 .lut_mask = 16'hFEFA;
defparam \Selector21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N20
cycloneive_lcell_comb \Selector21~8 (
// Equation(s):
// \Selector21~8_combout  = (\Selector21~7_combout ) # ((\Selector21~0_combout  & \Selector15~3_combout ))

	.dataa(gnd),
	.datab(\Selector21~0_combout ),
	.datac(\Selector15~3_combout ),
	.datad(\Selector21~7_combout ),
	.cin(gnd),
	.combout(\Selector21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~8 .lut_mask = 16'hFFC0;
defparam \Selector21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N24
cycloneive_lcell_comb \Selector20~1 (
// Equation(s):
// \Selector20~1_combout  = (\Selector20~0_combout  & ((\Selector15~3_combout ) # ((\ShiftRight0~30_combout  & \Selector23~0_combout )))) # (!\Selector20~0_combout  & (\ShiftRight0~30_combout  & (\Selector23~0_combout )))

	.dataa(\Selector20~0_combout ),
	.datab(\ShiftRight0~30_combout ),
	.datac(\Selector23~0_combout ),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~1 .lut_mask = 16'hEAC0;
defparam \Selector20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N2
cycloneive_lcell_comb \Selector20~4 (
// Equation(s):
// \Selector20~4_combout  = (!\input_b~63_combout  & (!\input_a~104_combout  & \Selector0~11_combout ))

	.dataa(gnd),
	.datab(input_b22),
	.datac(input_a20),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~4 .lut_mask = 16'h0300;
defparam \Selector20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N20
cycloneive_lcell_comb \Selector20~5 (
// Equation(s):
// \Selector20~5_combout  = (\Selector0~13_combout  & ((\Add1~22_combout ) # ((\Add0~22_combout  & \Selector0~12_combout )))) # (!\Selector0~13_combout  & (\Add0~22_combout  & (\Selector0~12_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Add0~22_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add1~22_combout ),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~5 .lut_mask = 16'hEAC0;
defparam \Selector20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N22
cycloneive_lcell_comb \Selector20~6 (
// Equation(s):
// \Selector20~6_combout  = (\Selector20~4_combout ) # ((\Selector20~5_combout ) # ((\Selector0~8_combout  & \input_a~104_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector20~4_combout ),
	.datac(input_a20),
	.datad(\Selector20~5_combout ),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~6 .lut_mask = 16'hFFEC;
defparam \Selector20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N18
cycloneive_lcell_comb \Selector20~2 (
// Equation(s):
// \Selector20~2_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~104_combout ))

	.dataa(gnd),
	.datab(\Selector0~9_combout ),
	.datac(input_a20),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~2 .lut_mask = 16'hFFC0;
defparam \Selector20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N4
cycloneive_lcell_comb \Selector20~3 (
// Equation(s):
// \Selector20~3_combout  = (\input_b~63_combout  & ((\Selector20~2_combout ) # ((!\input_a~104_combout  & \Selector0~10_combout )))) # (!\input_b~63_combout  & (((\input_a~104_combout  & \Selector0~10_combout ))))

	.dataa(input_b22),
	.datab(\Selector20~2_combout ),
	.datac(input_a20),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~3 .lut_mask = 16'hDA88;
defparam \Selector20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N0
cycloneive_lcell_comb \Selector20~7 (
// Equation(s):
// \Selector20~7_combout  = (\Selector20~6_combout ) # ((\Selector20~3_combout ) # ((\ShiftLeft0~82_combout  & \Selector16~9_combout )))

	.dataa(\Selector20~6_combout ),
	.datab(\Selector20~3_combout ),
	.datac(\ShiftLeft0~82_combout ),
	.datad(\Selector16~9_combout ),
	.cin(gnd),
	.combout(\Selector20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~7 .lut_mask = 16'hFEEE;
defparam \Selector20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N14
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (\Selector15~1_combout  & \ShiftRight0~70_combout )

	.dataa(gnd),
	.datab(\Selector15~1_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hCC00;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N22
cycloneive_lcell_comb \Selector9~6 (
// Equation(s):
// \Selector9~6_combout  = (\input_b~81_combout  & ((\ShiftLeft0~98_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~93_combout ))

	.dataa(\ShiftLeft0~93_combout ),
	.datab(input_b35),
	.datac(gnd),
	.datad(\ShiftLeft0~98_combout ),
	.cin(gnd),
	.combout(\Selector9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~6 .lut_mask = 16'hEE22;
defparam \Selector9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N4
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// \Selector9~1_combout  = (\Selector15~13_combout  & ((\input_b~81_combout  & (\ShiftLeft0~94_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~96_combout )))))

	.dataa(\ShiftLeft0~94_combout ),
	.datab(input_b35),
	.datac(\Selector15~13_combout ),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'hB080;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \Selector9~2 (
// Equation(s):
// \Selector9~2_combout  = (\input_b~33_combout  & (\Selector0~10_combout  & ((!\input_a~79_combout )))) # (!\input_b~33_combout  & ((\input_a~79_combout  & (\Selector0~10_combout )) # (!\input_a~79_combout  & ((\Selector0~11_combout )))))

	.dataa(input_b11),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~11_combout ),
	.datad(input_a9),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~2 .lut_mask = 16'h44D8;
defparam \Selector9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N22
cycloneive_lcell_comb \Selector9~3 (
// Equation(s):
// \Selector9~3_combout  = (\Selector0~13_combout  & ((\Add1~44_combout ) # ((\Selector0~12_combout  & Add01)))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & (Add01)))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(Add01),
	.datad(\Add1~44_combout ),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~3 .lut_mask = 16'hEAC0;
defparam \Selector9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N20
cycloneive_lcell_comb \Selector9~5 (
// Equation(s):
// \Selector9~5_combout  = (\Selector9~4_combout ) # ((\Selector9~2_combout ) # (\Selector9~3_combout ))

	.dataa(\Selector9~4_combout ),
	.datab(gnd),
	.datac(\Selector9~2_combout ),
	.datad(\Selector9~3_combout ),
	.cin(gnd),
	.combout(\Selector9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~5 .lut_mask = 16'hFFFA;
defparam \Selector9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N28
cycloneive_lcell_comb \Selector9~7 (
// Equation(s):
// \Selector9~7_combout  = (\Selector9~1_combout ) # ((\Selector9~5_combout ) # ((\Selector15~4_combout  & \Selector9~6_combout )))

	.dataa(\Selector15~4_combout ),
	.datab(\Selector9~6_combout ),
	.datac(\Selector9~1_combout ),
	.datad(\Selector9~5_combout ),
	.cin(gnd),
	.combout(\Selector9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~7 .lut_mask = 16'hFFF8;
defparam \Selector9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N18
cycloneive_lcell_comb \Selector8~3 (
// Equation(s):
// \Selector8~3_combout  = (\Selector0~12_combout  & ((Add02) # ((\Selector0~13_combout  & \Add1~46_combout )))) # (!\Selector0~12_combout  & (((\Selector0~13_combout  & \Add1~46_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(Add02),
	.datac(\Selector0~13_combout ),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\Selector8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~3 .lut_mask = 16'hF888;
defparam \Selector8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N8
cycloneive_lcell_comb \Selector8~4 (
// Equation(s):
// \Selector8~4_combout  = (\input_b~30_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~77_combout )))) # (!\input_b~30_combout  & (((\input_a~77_combout  & \Selector0~8_combout ))))

	.dataa(input_b10),
	.datab(\Selector0~9_combout ),
	.datac(input_a8),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~4 .lut_mask = 16'hFA80;
defparam \Selector8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N14
cycloneive_lcell_comb \Selector0~18 (
// Equation(s):
// \Selector0~18_combout  = (\input_b~81_combout  & ((\ShiftLeft0~84_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~79_combout ))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~18 .lut_mask = 16'hFA50;
defparam \Selector0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N18
cycloneive_lcell_comb \Selector8~9 (
// Equation(s):
// \Selector8~9_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & (\ShiftLeft0~80_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~83_combout )))))

	.dataa(input_b35),
	.datab(\ShiftLeft0~80_combout ),
	.datac(\Selector15~4_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\Selector8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~9 .lut_mask = 16'hD080;
defparam \Selector8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y29_N24
cycloneive_lcell_comb \Selector8~5 (
// Equation(s):
// \Selector8~5_combout  = (\input_b~30_combout  & (\Selector0~10_combout  & (!\input_a~77_combout ))) # (!\input_b~30_combout  & ((\input_a~77_combout  & (\Selector0~10_combout )) # (!\input_a~77_combout  & ((\Selector0~11_combout )))))

	.dataa(input_b10),
	.datab(\Selector0~10_combout ),
	.datac(input_a8),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~5 .lut_mask = 16'h4D48;
defparam \Selector8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N30
cycloneive_lcell_comb \Selector8~6 (
// Equation(s):
// \Selector8~6_combout  = (\Selector8~9_combout ) # ((\Selector8~5_combout ) # ((\Selector15~1_combout  & \ShiftRight0~73_combout )))

	.dataa(\Selector15~1_combout ),
	.datab(\Selector8~9_combout ),
	.datac(\Selector8~5_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\Selector8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~6 .lut_mask = 16'hFEFC;
defparam \Selector8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N14
cycloneive_lcell_comb \Selector8~7 (
// Equation(s):
// \Selector8~7_combout  = (\Selector8~4_combout ) # ((\Selector8~6_combout ) # ((\Selector15~13_combout  & \Selector0~18_combout )))

	.dataa(\Selector8~4_combout ),
	.datab(\Selector15~13_combout ),
	.datac(\Selector0~18_combout ),
	.datad(\Selector8~6_combout ),
	.cin(gnd),
	.combout(\Selector8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~7 .lut_mask = 16'hFFEA;
defparam \Selector8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N12
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (\input_b~81_combout  & ((\ShiftLeft0~70_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~62_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftLeft0~62_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N14
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (!\ShiftLeft0~104_combout  & (\Selector15~6_combout  & (!\input_b~79_combout  & \ShiftLeft0~21_combout )))

	.dataa(\ShiftLeft0~104_combout ),
	.datab(\Selector15~6_combout ),
	.datac(input_b33),
	.datad(\ShiftLeft0~21_combout ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'h0400;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N16
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & ((\ShiftLeft0~49_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~52_combout ))))

	.dataa(\ShiftLeft0~52_combout ),
	.datab(input_b35),
	.datac(\Selector15~4_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'hE020;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N8
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// \Selector14~2_combout  = (\input_a~89_combout  & (((!\input_b~48_combout  & \Selector0~10_combout )))) # (!\input_a~89_combout  & ((\input_b~48_combout  & ((\Selector0~10_combout ))) # (!\input_b~48_combout  & (\Selector0~11_combout ))))

	.dataa(input_a14),
	.datab(\Selector0~11_combout ),
	.datac(input_b16),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'h5E04;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N10
cycloneive_lcell_comb \Selector14~3 (
// Equation(s):
// \Selector14~3_combout  = (\Add1~34_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add0~34_combout )))) # (!\Add1~34_combout  & (((\Selector0~12_combout  & \Add0~34_combout ))))

	.dataa(\Add1~34_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add0~34_combout ),
	.cin(gnd),
	.combout(\Selector14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~3 .lut_mask = 16'hF888;
defparam \Selector14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N24
cycloneive_lcell_comb \Selector14~4 (
// Equation(s):
// \Selector14~4_combout  = (\input_a~89_combout  & ((\Selector0~8_combout ) # ((\input_b~48_combout  & \Selector0~9_combout )))) # (!\input_a~89_combout  & (\input_b~48_combout  & ((\Selector0~8_combout ))))

	.dataa(input_a14),
	.datab(input_b16),
	.datac(\Selector0~9_combout ),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~4 .lut_mask = 16'hEE80;
defparam \Selector14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N18
cycloneive_lcell_comb \Selector14~5 (
// Equation(s):
// \Selector14~5_combout  = (\Selector14~2_combout ) # ((\Selector14~3_combout ) # (\Selector14~4_combout ))

	.dataa(gnd),
	.datab(\Selector14~2_combout ),
	.datac(\Selector14~3_combout ),
	.datad(\Selector14~4_combout ),
	.cin(gnd),
	.combout(\Selector14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~5 .lut_mask = 16'hFFFC;
defparam \Selector14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N26
cycloneive_lcell_comb \Selector14~6 (
// Equation(s):
// \Selector14~6_combout  = (\Selector14~1_combout ) # ((\Selector14~5_combout ) # ((\ShiftRight0~27_combout  & \Selector15~1_combout )))

	.dataa(\ShiftRight0~27_combout ),
	.datab(\Selector14~1_combout ),
	.datac(\Selector15~1_combout ),
	.datad(\Selector14~5_combout ),
	.cin(gnd),
	.combout(\Selector14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~6 .lut_mask = 16'hFFEC;
defparam \Selector14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N30
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (\input_b~83_combout  & (\ShiftLeft0~31_combout )) # (!\input_b~83_combout  & ((\ShiftLeft0~33_combout )))

	.dataa(input_b37),
	.datab(gnd),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N8
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\input_b~83_combout  & ((\ShiftLeft0~45_combout ))) # (!\input_b~83_combout  & (\ShiftLeft0~30_combout ))

	.dataa(input_b37),
	.datab(\ShiftLeft0~30_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y27_N12
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (\input_b~81_combout  & ((\ShiftLeft0~93_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~94_combout ))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftLeft0~94_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N4
cycloneive_lcell_comb \Selector13~0 (
// Equation(s):
// \Selector13~0_combout  = (\ShiftLeft0~73_combout  & (\Selector15~6_combout  & \ShiftLeft0~103_combout ))

	.dataa(\ShiftLeft0~73_combout ),
	.datab(\Selector15~6_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~0 .lut_mask = 16'h8800;
defparam \Selector13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N0
cycloneive_lcell_comb \Selector13~1 (
// Equation(s):
// \Selector13~1_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & (\ShiftLeft0~74_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~98_combout )))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(\Selector15~4_combout ),
	.datac(input_b35),
	.datad(\ShiftLeft0~98_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~1 .lut_mask = 16'h8C80;
defparam \Selector13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N26
cycloneive_lcell_comb \Selector13~4 (
// Equation(s):
// \Selector13~4_combout  = (\input_b~45_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_a~87_combout )))) # (!\input_b~45_combout  & (((\Selector0~8_combout  & \input_a~87_combout ))))

	.dataa(input_b15),
	.datab(\Selector0~9_combout ),
	.datac(\Selector0~8_combout ),
	.datad(input_a13),
	.cin(gnd),
	.combout(\Selector13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~4 .lut_mask = 16'hF8A0;
defparam \Selector13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N12
cycloneive_lcell_comb \Selector13~3 (
// Equation(s):
// \Selector13~3_combout  = (\Add1~36_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add0~36_combout )))) # (!\Add1~36_combout  & (((\Selector0~12_combout  & \Add0~36_combout ))))

	.dataa(\Add1~36_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add0~36_combout ),
	.cin(gnd),
	.combout(\Selector13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~3 .lut_mask = 16'hF888;
defparam \Selector13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N20
cycloneive_lcell_comb \Selector13~5 (
// Equation(s):
// \Selector13~5_combout  = (\Selector13~2_combout ) # ((\Selector13~4_combout ) # (\Selector13~3_combout ))

	.dataa(\Selector13~2_combout ),
	.datab(gnd),
	.datac(\Selector13~4_combout ),
	.datad(\Selector13~3_combout ),
	.cin(gnd),
	.combout(\Selector13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~5 .lut_mask = 16'hFFFA;
defparam \Selector13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N2
cycloneive_lcell_comb \Selector13~6 (
// Equation(s):
// \Selector13~6_combout  = (\Selector13~1_combout ) # ((\Selector13~5_combout ) # ((\ShiftRight0~79_combout  & \Selector15~1_combout )))

	.dataa(\Selector13~1_combout ),
	.datab(\Selector13~5_combout ),
	.datac(\ShiftRight0~79_combout ),
	.datad(\Selector15~1_combout ),
	.cin(gnd),
	.combout(\Selector13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~6 .lut_mask = 16'hFEEE;
defparam \Selector13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N12
cycloneive_lcell_comb \Selector12~0 (
// Equation(s):
// \Selector12~0_combout  = (\ShiftLeft0~103_combout  & (\ShiftLeft0~23_combout  & \Selector15~6_combout ))

	.dataa(\ShiftLeft0~103_combout ),
	.datab(\ShiftLeft0~23_combout ),
	.datac(gnd),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~0 .lut_mask = 16'h8800;
defparam \Selector12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N18
cycloneive_lcell_comb \Selector12~2 (
// Equation(s):
// \Selector12~2_combout  = (\input_a~85_combout  & (!\input_b~42_combout  & ((\Selector0~10_combout )))) # (!\input_a~85_combout  & ((\input_b~42_combout  & ((\Selector0~10_combout ))) # (!\input_b~42_combout  & (\Selector0~11_combout ))))

	.dataa(input_a12),
	.datab(input_b14),
	.datac(\Selector0~11_combout ),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~2 .lut_mask = 16'h7610;
defparam \Selector12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N14
cycloneive_lcell_comb \Selector12~4 (
// Equation(s):
// \Selector12~4_combout  = (\Selector0~8_combout  & ((\input_b~42_combout ) # ((\input_a~85_combout )))) # (!\Selector0~8_combout  & (\input_b~42_combout  & (\Selector0~9_combout  & \input_a~85_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(input_b14),
	.datac(\Selector0~9_combout ),
	.datad(input_a12),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~4 .lut_mask = 16'hEA88;
defparam \Selector12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N16
cycloneive_lcell_comb \Selector12~3 (
// Equation(s):
// \Selector12~3_combout  = (\Add0~38_combout  & ((\Selector0~12_combout ) # ((\Selector0~13_combout  & \Add1~38_combout )))) # (!\Add0~38_combout  & (\Selector0~13_combout  & ((\Add1~38_combout ))))

	.dataa(\Add0~38_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~3 .lut_mask = 16'hECA0;
defparam \Selector12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N28
cycloneive_lcell_comb \Selector12~5 (
// Equation(s):
// \Selector12~5_combout  = (\Selector12~2_combout ) # ((\Selector12~4_combout ) # (\Selector12~3_combout ))

	.dataa(gnd),
	.datab(\Selector12~2_combout ),
	.datac(\Selector12~4_combout ),
	.datad(\Selector12~3_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~5 .lut_mask = 16'hFFFC;
defparam \Selector12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y28_N18
cycloneive_lcell_comb \Selector12~1 (
// Equation(s):
// \Selector12~1_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & (\ShiftLeft0~76_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~80_combout )))))

	.dataa(\ShiftLeft0~76_combout ),
	.datab(\ShiftLeft0~80_combout ),
	.datac(\Selector15~4_combout ),
	.datad(input_b35),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~1 .lut_mask = 16'hA0C0;
defparam \Selector12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y28_N28
cycloneive_lcell_comb \Selector12~6 (
// Equation(s):
// \Selector12~6_combout  = (\Selector12~5_combout ) # ((\Selector12~1_combout ) # ((\ShiftLeft0~85_combout  & \Selector15~13_combout )))

	.dataa(\ShiftLeft0~85_combout ),
	.datab(\Selector15~13_combout ),
	.datac(\Selector12~5_combout ),
	.datad(\Selector12~1_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~6 .lut_mask = 16'hFFF8;
defparam \Selector12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y26_N18
cycloneive_lcell_comb \Selector23~2 (
// Equation(s):
// \Selector23~2_combout  = (\ShiftLeft0~91_combout  & \Selector16~9_combout )

	.dataa(\ShiftLeft0~91_combout ),
	.datab(gnd),
	.datac(\Selector16~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~2 .lut_mask = 16'hA0A0;
defparam \Selector23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y27_N16
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\input_b~85_combout  & (\input_a~85_combout )) # (!\input_b~85_combout  & ((\input_a~87_combout )))

	.dataa(input_a12),
	.datab(input_b39),
	.datac(gnd),
	.datad(input_a13),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hBB88;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N30
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\input_b~83_combout  & (\ShiftRight0~41_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~42_combout )))

	.dataa(gnd),
	.datab(input_b37),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N10
cycloneive_lcell_comb \Selector23~1 (
// Equation(s):
// \Selector23~1_combout  = (\input_b~81_combout  & ((\ShiftRight0~59_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~43_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~59_combout ),
	.cin(gnd),
	.combout(\Selector23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~1 .lut_mask = 16'hFC30;
defparam \Selector23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N24
cycloneive_lcell_comb \Selector23~5 (
// Equation(s):
// \Selector23~5_combout  = (\Selector0~11_combout  & (!\input_a~113_combout  & !\input_b~69_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(input_a23),
	.datac(input_b25),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~5 .lut_mask = 16'h0202;
defparam \Selector23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N2
cycloneive_lcell_comb \Selector23~6 (
// Equation(s):
// \Selector23~6_combout  = (\Selector0~12_combout  & ((\Add0~16_combout ) # ((\Add1~16_combout  & \Selector0~13_combout )))) # (!\Selector0~12_combout  & (\Add1~16_combout  & (\Selector0~13_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add1~16_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Add0~16_combout ),
	.cin(gnd),
	.combout(\Selector23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~6 .lut_mask = 16'hEAC0;
defparam \Selector23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N4
cycloneive_lcell_comb \Selector23~7 (
// Equation(s):
// \Selector23~7_combout  = (\Selector23~5_combout ) # ((\Selector23~6_combout ) # ((\Selector0~8_combout  & \input_a~113_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector23~5_combout ),
	.datac(input_a23),
	.datad(\Selector23~6_combout ),
	.cin(gnd),
	.combout(\Selector23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~7 .lut_mask = 16'hFFEC;
defparam \Selector23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y28_N22
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\input_b~83_combout  & (\ShiftRight0~48_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~49_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~48_combout ),
	.datac(input_b37),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N20
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\input_b~83_combout  & (\ShiftRight0~44_combout )) # (!\input_b~83_combout  & ((\ShiftRight0~45_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~44_combout ),
	.datac(\ShiftRight0~45_combout ),
	.datad(input_b37),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N30
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\input_b~81_combout  & ((\ShiftRight0~46_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~50_combout ))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftRight0~50_combout ),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hFC30;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N22
cycloneive_lcell_comb \Selector23~8 (
// Equation(s):
// \Selector23~8_combout  = (\Selector23~4_combout ) # ((\Selector23~7_combout ) # ((\Selector16~0_combout  & \ShiftRight0~85_combout )))

	.dataa(\Selector23~4_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector23~7_combout ),
	.datad(\ShiftRight0~85_combout ),
	.cin(gnd),
	.combout(\Selector23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~8 .lut_mask = 16'hFEFA;
defparam \Selector23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y26_N28
cycloneive_lcell_comb \Selector23~9 (
// Equation(s):
// \Selector23~9_combout  = (\Selector23~8_combout ) # ((\Selector23~1_combout  & \Selector15~3_combout ))

	.dataa(\Selector23~1_combout ),
	.datab(gnd),
	.datac(\Selector23~8_combout ),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~9 .lut_mask = 16'hFAF0;
defparam \Selector23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N4
cycloneive_lcell_comb \Selector19~7 (
// Equation(s):
// \Selector19~7_combout  = (ALUOP_ID_0 & (\input_b~77_combout  & (\ShiftLeft0~103_combout  & \Selector15~0_combout )))

	.dataa(ALUOP_ID_0),
	.datab(input_b31),
	.datac(\ShiftLeft0~103_combout ),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~7 .lut_mask = 16'h8000;
defparam \Selector19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N26
cycloneive_lcell_comb \Selector19~0 (
// Equation(s):
// \Selector19~0_combout  = (\Selector15~3_combout  & ((\input_b~81_combout  & (\ShiftRight0~56_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~59_combout )))))

	.dataa(\ShiftRight0~56_combout ),
	.datab(input_b35),
	.datac(\Selector15~3_combout ),
	.datad(\ShiftRight0~59_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~0 .lut_mask = 16'hB080;
defparam \Selector19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N18
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\input_b~81_combout  & (\ShiftRight0~43_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~46_combout )))

	.dataa(input_b35),
	.datab(gnd),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N8
cycloneive_lcell_comb \Selector19~1 (
// Equation(s):
// \Selector19~1_combout  = (\input_b~61_combout  & ((\Selector0~8_combout ) # ((\input_a~101_combout  & \Selector0~9_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(input_a19),
	.datac(\Selector0~9_combout ),
	.datad(input_b21),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~1 .lut_mask = 16'hEA00;
defparam \Selector19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N26
cycloneive_lcell_comb \Selector19~2 (
// Equation(s):
// \Selector19~2_combout  = (\Selector19~1_combout ) # ((\Selector0~10_combout  & (\input_b~61_combout  $ (\input_a~101_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(input_b21),
	.datac(\Selector19~1_combout ),
	.datad(input_a19),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~2 .lut_mask = 16'hF2F8;
defparam \Selector19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N22
cycloneive_lcell_comb \Selector19~6 (
// Equation(s):
// \Selector19~6_combout  = (\Selector19~5_combout ) # ((\Selector19~2_combout ) # ((\ShiftRight0~47_combout  & \Selector16~0_combout )))

	.dataa(\Selector19~5_combout ),
	.datab(\ShiftRight0~47_combout ),
	.datac(\Selector19~2_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~6 .lut_mask = 16'hFEFA;
defparam \Selector19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N18
cycloneive_lcell_comb \Selector19~8 (
// Equation(s):
// \Selector19~8_combout  = (\Selector19~0_combout ) # ((\Selector19~6_combout ) # ((\ShiftRight0~40_combout  & \Selector19~7_combout )))

	.dataa(\ShiftRight0~40_combout ),
	.datab(\Selector19~7_combout ),
	.datac(\Selector19~0_combout ),
	.datad(\Selector19~6_combout ),
	.cin(gnd),
	.combout(\Selector19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~8 .lut_mask = 16'hFFF8;
defparam \Selector19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y27_N22
cycloneive_lcell_comb \Selector10~2 (
// Equation(s):
// \Selector10~2_combout  = (\input_b~81_combout  & (\ShiftLeft0~52_combout )) # (!\input_b~81_combout  & ((\ShiftLeft0~70_combout )))

	.dataa(gnd),
	.datab(input_b35),
	.datac(\ShiftLeft0~52_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~2 .lut_mask = 16'hF3C0;
defparam \Selector10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N10
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\input_b~79_combout  & (\ShiftLeft0~67_combout )) # (!\input_b~79_combout  & ((\Selector10~2_combout )))

	.dataa(input_b33),
	.datab(gnd),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\Selector10~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \Selector18~4 (
// Equation(s):
// \Selector18~4_combout  = (\Add1~26_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add0~26_combout )))) # (!\Add1~26_combout  & (\Selector0~12_combout  & ((\Add0~26_combout ))))

	.dataa(\Add1~26_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Add0~26_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~4 .lut_mask = 16'hECA0;
defparam \Selector18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \Selector18~3 (
// Equation(s):
// \Selector18~3_combout  = (!\input_b~59_combout  & (!\input_a~98_combout  & \Selector0~11_combout ))

	.dataa(input_b20),
	.datab(input_a18),
	.datac(gnd),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~3 .lut_mask = 16'h1100;
defparam \Selector18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \Selector18~5 (
// Equation(s):
// \Selector18~5_combout  = (\Selector18~4_combout ) # ((\Selector18~3_combout ) # ((\Selector0~8_combout  & \input_a~98_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(input_a18),
	.datac(\Selector18~4_combout ),
	.datad(\Selector18~3_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~5 .lut_mask = 16'hFFF8;
defparam \Selector18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \Selector18~6 (
// Equation(s):
// \Selector18~6_combout  = (\Selector18~2_combout ) # ((\Selector18~5_combout ) # ((\ShiftRight0~74_combout  & \Selector16~0_combout )))

	.dataa(\Selector18~2_combout ),
	.datab(\Selector18~5_combout ),
	.datac(\ShiftRight0~74_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~6 .lut_mask = 16'hFEEE;
defparam \Selector18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N6
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// \Selector18~0_combout  = (\Selector15~3_combout  & ((\input_b~81_combout  & (\ShiftRight0~19_combout )) # (!\input_b~81_combout  & ((\ShiftRight0~23_combout )))))

	.dataa(\ShiftRight0~19_combout ),
	.datab(input_b35),
	.datac(\Selector15~3_combout ),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'hB080;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N28
cycloneive_lcell_comb \Selector18~7 (
// Equation(s):
// \Selector18~7_combout  = (\Selector18~6_combout ) # ((\Selector18~0_combout ) # ((\ShiftRight0~16_combout  & \Selector19~7_combout )))

	.dataa(\ShiftRight0~16_combout ),
	.datab(\Selector19~7_combout ),
	.datac(\Selector18~6_combout ),
	.datad(\Selector18~0_combout ),
	.cin(gnd),
	.combout(\Selector18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~7 .lut_mask = 16'hFFF8;
defparam \Selector18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y27_N10
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (\input_b~79_combout  & (\ShiftLeft0~75_combout )) # (!\input_b~79_combout  & ((\Selector9~6_combout )))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(gnd),
	.datac(input_b33),
	.datad(\Selector9~6_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N8
cycloneive_lcell_comb \Selector17~0 (
// Equation(s):
// \Selector17~0_combout  = (\ShiftRight0~38_combout  & (!\ShiftLeft0~104_combout  & \Selector23~0_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~38_combout ),
	.datac(\ShiftLeft0~104_combout ),
	.datad(\Selector23~0_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~0 .lut_mask = 16'h0C00;
defparam \Selector17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N20
cycloneive_lcell_comb \Selector17~4 (
// Equation(s):
// \Selector17~4_combout  = (\input_a~95_combout  & ((\Selector0~8_combout ) # ((\input_b~57_combout  & \Selector0~9_combout )))) # (!\input_a~95_combout  & (\Selector0~8_combout  & (\input_b~57_combout )))

	.dataa(input_a17),
	.datab(\Selector0~8_combout ),
	.datac(input_b19),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~4 .lut_mask = 16'hE8C8;
defparam \Selector17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N6
cycloneive_lcell_comb \Selector17~2 (
// Equation(s):
// \Selector17~2_combout  = (\input_b~57_combout  & (\Selector0~10_combout  & ((!\input_a~95_combout )))) # (!\input_b~57_combout  & ((\input_a~95_combout  & (\Selector0~10_combout )) # (!\input_a~95_combout  & ((\Selector0~11_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(input_b19),
	.datac(\Selector0~11_combout ),
	.datad(input_a17),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~2 .lut_mask = 16'h22B8;
defparam \Selector17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N4
cycloneive_lcell_comb \Selector17~5 (
// Equation(s):
// \Selector17~5_combout  = (\Selector17~3_combout ) # ((\Selector17~4_combout ) # (\Selector17~2_combout ))

	.dataa(\Selector17~3_combout ),
	.datab(gnd),
	.datac(\Selector17~4_combout ),
	.datad(\Selector17~2_combout ),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~5 .lut_mask = 16'hFFFA;
defparam \Selector17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N12
cycloneive_lcell_comb \Selector17~1 (
// Equation(s):
// \Selector17~1_combout  = (\Selector15~3_combout  & ((\input_b~81_combout  & ((\ShiftRight0~67_combout ))) # (!\input_b~81_combout  & (\ShiftRight0~68_combout ))))

	.dataa(\ShiftRight0~68_combout ),
	.datab(input_b35),
	.datac(\ShiftRight0~67_combout ),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~1 .lut_mask = 16'hE200;
defparam \Selector17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N26
cycloneive_lcell_comb \Selector17~6 (
// Equation(s):
// \Selector17~6_combout  = (\Selector17~5_combout ) # ((\Selector17~1_combout ) # ((\ShiftRight0~65_combout  & \Selector16~0_combout )))

	.dataa(\Selector17~5_combout ),
	.datab(\ShiftRight0~65_combout ),
	.datac(\Selector16~0_combout ),
	.datad(\Selector17~1_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~6 .lut_mask = 16'hFFEA;
defparam \Selector17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N2
cycloneive_lcell_comb \Selector0~27 (
// Equation(s):
// \Selector0~27_combout  = (Add1 & \Selector0~13_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Add1),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~27 .lut_mask = 16'hF000;
defparam \Selector0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N24
cycloneive_lcell_comb \Selector0~20 (
// Equation(s):
// \Selector0~20_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & \input_b~6_combout ))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(gnd),
	.datad(input_b2),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~20 .lut_mask = 16'hEEAA;
defparam \Selector0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N22
cycloneive_lcell_comb \Selector0~21 (
// Equation(s):
// \Selector0~21_combout  = (\input_a~61_combout  & ((\Selector0~20_combout ) # ((!\ShiftLeft0~87_combout  & \Selector15~1_combout ))))

	.dataa(input_a),
	.datab(\ShiftLeft0~87_combout ),
	.datac(\Selector15~1_combout ),
	.datad(\Selector0~20_combout ),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~21 .lut_mask = 16'hAA20;
defparam \Selector0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N2
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (\input_b~81_combout ) # ((\input_b~85_combout  & !\input_b~83_combout ))

	.dataa(gnd),
	.datab(input_b39),
	.datac(input_b37),
	.datad(input_b35),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'hFF0C;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N20
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\input_b~85_combout  & (\input_a~67_combout )) # (!\input_b~85_combout  & ((\input_a~65_combout )))

	.dataa(input_a3),
	.datab(input_a2),
	.datac(input_b39),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hACAC;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N16
cycloneive_lcell_comb \Selector0~22 (
// Equation(s):
// \Selector0~22_combout  = (\ShiftLeft0~104_combout  & ((\ShiftLeft0~59_combout ) # ((\Selector1~1_combout )))) # (!\ShiftLeft0~104_combout  & (((\input_a~61_combout  & !\Selector1~1_combout ))))

	.dataa(\ShiftLeft0~104_combout ),
	.datab(\ShiftLeft0~59_combout ),
	.datac(input_a),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~22 .lut_mask = 16'hAAD8;
defparam \Selector0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N6
cycloneive_lcell_comb \Selector0~23 (
// Equation(s):
// \Selector0~23_combout  = (\Selector1~1_combout  & ((\Selector0~22_combout  & (\ShiftLeft0~86_combout )) # (!\Selector0~22_combout  & ((\input_a~63_combout ))))) # (!\Selector1~1_combout  & (((\Selector0~22_combout ))))

	.dataa(\ShiftLeft0~86_combout ),
	.datab(input_a1),
	.datac(\Selector1~1_combout ),
	.datad(\Selector0~22_combout ),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~23 .lut_mask = 16'hAFC0;
defparam \Selector0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N8
cycloneive_lcell_comb \Selector0~24 (
// Equation(s):
// \Selector0~24_combout  = (\ShiftLeft0~88_combout  & ((\Selector15~6_combout ) # ((\Selector15~13_combout  & \Selector0~23_combout )))) # (!\ShiftLeft0~88_combout  & (\Selector15~13_combout  & (\Selector0~23_combout )))

	.dataa(\ShiftLeft0~88_combout ),
	.datab(\Selector15~13_combout ),
	.datac(\Selector0~23_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~24 .lut_mask = 16'hEAC0;
defparam \Selector0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N30
cycloneive_lcell_comb \Selector0~19 (
// Equation(s):
// \Selector0~19_combout  = (\input_a~61_combout  & (\Selector0~10_combout  & ((!\input_b~6_combout )))) # (!\input_a~61_combout  & ((\input_b~6_combout  & (\Selector0~10_combout )) # (!\input_b~6_combout  & ((\Selector0~11_combout )))))

	.dataa(input_a),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~11_combout ),
	.datad(input_b2),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~19 .lut_mask = 16'h44D8;
defparam \Selector0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N2
cycloneive_lcell_comb \Selector0~25 (
// Equation(s):
// \Selector0~25_combout  = (\Selector0~8_combout  & ((\input_b~6_combout ) # ((\Selector0~18_combout  & \Selector15~4_combout )))) # (!\Selector0~8_combout  & (\Selector0~18_combout  & ((\Selector15~4_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~18_combout ),
	.datac(input_b2),
	.datad(\Selector15~4_combout ),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~25 .lut_mask = 16'hECA0;
defparam \Selector0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N0
cycloneive_lcell_comb \Selector0~26 (
// Equation(s):
// \Selector0~26_combout  = (\Selector0~21_combout ) # ((\Selector0~24_combout ) # ((\Selector0~19_combout ) # (\Selector0~25_combout )))

	.dataa(\Selector0~21_combout ),
	.datab(\Selector0~24_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Selector0~25_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~26 .lut_mask = 16'hFFFE;
defparam \Selector0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y30_N22
cycloneive_lcell_comb \Selector1~6 (
// Equation(s):
// \Selector1~6_combout  = (\Selector1~5_combout  & (((\ShiftLeft0~97_combout ) # (!\Selector1~1_combout )))) # (!\Selector1~5_combout  & (\input_a~65_combout  & (\Selector1~1_combout )))

	.dataa(\Selector1~5_combout ),
	.datab(input_a2),
	.datac(\Selector1~1_combout ),
	.datad(\ShiftLeft0~97_combout ),
	.cin(gnd),
	.combout(\Selector1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~6 .lut_mask = 16'hEA4A;
defparam \Selector1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N12
cycloneive_lcell_comb \Selector1~7 (
// Equation(s):
// \Selector1~7_combout  = (\ShiftLeft0~101_combout  & ((\Selector15~6_combout ) # ((\Selector15~13_combout  & \Selector1~6_combout )))) # (!\ShiftLeft0~101_combout  & (\Selector15~13_combout  & (\Selector1~6_combout )))

	.dataa(\ShiftLeft0~101_combout ),
	.datab(\Selector15~13_combout ),
	.datac(\Selector1~6_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~7 .lut_mask = 16'hEAC0;
defparam \Selector1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N16
cycloneive_lcell_comb \Selector1~3 (
// Equation(s):
// \Selector1~3_combout  = (\Selector0~8_combout  & ((\input_a~63_combout ) # ((\input_b~9_combout )))) # (!\Selector0~8_combout  & (\input_a~63_combout  & (\Selector0~9_combout  & \input_b~9_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(input_a1),
	.datac(\Selector0~9_combout ),
	.datad(input_b3),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~3 .lut_mask = 16'hEA88;
defparam \Selector1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N26
cycloneive_lcell_comb \Selector1~2 (
// Equation(s):
// \Selector1~2_combout  = (\input_b~9_combout  & (((!\input_a~63_combout  & \Selector0~10_combout )))) # (!\input_b~9_combout  & ((\input_a~63_combout  & ((\Selector0~10_combout ))) # (!\input_a~63_combout  & (\Selector0~11_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(input_b3),
	.datac(input_a1),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~2 .lut_mask = 16'h3E02;
defparam \Selector1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N6
cycloneive_lcell_comb \Selector1~4 (
// Equation(s):
// \Selector1~4_combout  = (\Selector15~4_combout  & ((\input_b~81_combout  & ((\ShiftLeft0~94_combout ))) # (!\input_b~81_combout  & (\ShiftLeft0~96_combout ))))

	.dataa(input_b35),
	.datab(\ShiftLeft0~96_combout ),
	.datac(\ShiftLeft0~94_combout ),
	.datad(\Selector15~4_combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~4 .lut_mask = 16'hE400;
defparam \Selector1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y29_N10
cycloneive_lcell_comb \Selector1~8 (
// Equation(s):
// \Selector1~8_combout  = (\Selector1~7_combout ) # ((\Selector1~3_combout ) # ((\Selector1~2_combout ) # (\Selector1~4_combout )))

	.dataa(\Selector1~7_combout ),
	.datab(\Selector1~3_combout ),
	.datac(\Selector1~2_combout ),
	.datad(\Selector1~4_combout ),
	.cin(gnd),
	.combout(\Selector1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~8 .lut_mask = 16'hFFFE;
defparam \Selector1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N26
cycloneive_lcell_comb \Selector1~9 (
// Equation(s):
// \Selector1~9_combout  = (\Selector15~1_combout  & (!\input_b~79_combout  & (!\ShiftLeft0~104_combout  & \ShiftRight0~38_combout )))

	.dataa(\Selector15~1_combout ),
	.datab(input_b33),
	.datac(\ShiftLeft0~104_combout ),
	.datad(\ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\Selector1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~9 .lut_mask = 16'h0200;
defparam \Selector1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N16
cycloneive_lcell_comb \Selector1~10 (
// Equation(s):
// \Selector1~10_combout  = (\Selector1~9_combout ) # ((\Selector0~13_combout  & \Add1~60_combout ))

	.dataa(gnd),
	.datab(\Selector0~13_combout ),
	.datac(\Selector1~9_combout ),
	.datad(\Add1~60_combout ),
	.cin(gnd),
	.combout(\Selector1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~10 .lut_mask = 16'hFCF0;
defparam \Selector1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N20
cycloneive_lcell_comb \Equal11~10 (
// Equation(s):
// \Equal11~10_combout  = (!Selector1 & !Selector0)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector1),
	.datad(Selector0),
	.cin(gnd),
	.combout(\Equal11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~10 .lut_mask = 16'h000F;
defparam \Equal11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \Equal11~7 (
// Equation(s):
// \Equal11~7_combout  = (!Selector23 & (!Selector17 & (!Selector18 & !Selector19)))

	.dataa(Selector23),
	.datab(Selector17),
	.datac(Selector18),
	.datad(Selector19),
	.cin(gnd),
	.combout(\Equal11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~7 .lut_mask = 16'h0001;
defparam \Equal11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \Equal11~8 (
// Equation(s):
// \Equal11~8_combout  = (!Selector13 & (!Selector14 & (!Selector12 & \Equal11~7_combout )))

	.dataa(Selector13),
	.datab(Selector14),
	.datac(Selector12),
	.datad(\Equal11~7_combout ),
	.cin(gnd),
	.combout(\Equal11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~8 .lut_mask = 16'h0100;
defparam \Equal11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \Equal11~6 (
// Equation(s):
// \Equal11~6_combout  = (!Selector21 & (!Selector20 & (!Selector11 & !Selector10)))

	.dataa(Selector21),
	.datab(Selector20),
	.datac(Selector11),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Equal11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~6 .lut_mask = 16'h0001;
defparam \Equal11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N8
cycloneive_lcell_comb \Equal11~9 (
// Equation(s):
// \Equal11~9_combout  = (!Selector8 & (!Selector9 & (\Equal11~8_combout  & \Equal11~6_combout )))

	.dataa(Selector8),
	.datab(Selector9),
	.datac(\Equal11~8_combout ),
	.datad(\Equal11~6_combout ),
	.cin(gnd),
	.combout(\Equal11~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~9 .lut_mask = 16'h1000;
defparam \Equal11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N18
cycloneive_lcell_comb \Equal11~3 (
// Equation(s):
// \Equal11~3_combout  = (Selector15) # ((Selector29) # (Selector5))

	.dataa(gnd),
	.datab(Selector15),
	.datac(Selector29),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Equal11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~3 .lut_mask = 16'hFFFC;
defparam \Equal11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N8
cycloneive_lcell_comb \Equal11~2 (
// Equation(s):
// \Equal11~2_combout  = (!Selector7 & (!Selector16 & !Selector6))

	.dataa(gnd),
	.datab(Selector7),
	.datac(Selector16),
	.datad(Selector6),
	.cin(gnd),
	.combout(\Equal11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~2 .lut_mask = 16'h0003;
defparam \Equal11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N24
cycloneive_lcell_comb \Equal11~1 (
// Equation(s):
// \Equal11~1_combout  = (!Selector26 & (!Selector27 & (!Selector25 & !Selector24)))

	.dataa(Selector26),
	.datab(Selector27),
	.datac(Selector25),
	.datad(Selector24),
	.cin(gnd),
	.combout(\Equal11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~1 .lut_mask = 16'h0001;
defparam \Equal11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N4
cycloneive_lcell_comb \Equal11~4 (
// Equation(s):
// \Equal11~4_combout  = (!Selector4 & (!\Equal11~3_combout  & (\Equal11~2_combout  & \Equal11~1_combout )))

	.dataa(Selector4),
	.datab(\Equal11~3_combout ),
	.datac(\Equal11~2_combout ),
	.datad(\Equal11~1_combout ),
	.cin(gnd),
	.combout(\Equal11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~4 .lut_mask = 16'h1000;
defparam \Equal11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N10
cycloneive_lcell_comb \Equal11~0 (
// Equation(s):
// \Equal11~0_combout  = (!Selector30 & (!Selector22 & !Selector2))

	.dataa(gnd),
	.datab(Selector30),
	.datac(Selector22),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Equal11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~0 .lut_mask = 16'h0003;
defparam \Equal11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N30
cycloneive_lcell_comb \Equal11~5 (
// Equation(s):
// \Equal11~5_combout  = (!Selector3 & (!Selector28 & (\Equal11~4_combout  & \Equal11~0_combout )))

	.dataa(Selector3),
	.datab(Selector28),
	.datac(\Equal11~4_combout ),
	.datad(\Equal11~0_combout ),
	.cin(gnd),
	.combout(\Equal11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~5 .lut_mask = 16'h1000;
defparam \Equal11~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	Instr_IF_30,
	Instr_IF_28,
	Instr_IF_26,
	Instr_IF_27,
	Selector14,
	Instr_IF_29,
	Instr_IF_5,
	Instr_IF_4,
	Instr_IF_2,
	Instr_IF_3,
	Instr_IF_0,
	Selector11,
	Instr_IF_1,
	WideOr4,
	WideOr41,
	Instr_IF_31,
	input_hazard_Reg_ID,
	WideOr21,
	Selector141,
	WideOr211,
	WideOr212,
	WideOr14,
	WideOr6,
	WideOr61,
	WideOr33,
	Decoder0,
	WideOr11,
	devpor,
	devclrn,
	devoe);
input 	Instr_IF_30;
input 	Instr_IF_28;
input 	Instr_IF_26;
input 	Instr_IF_27;
output 	Selector14;
input 	Instr_IF_29;
input 	Instr_IF_5;
input 	Instr_IF_4;
input 	Instr_IF_2;
input 	Instr_IF_3;
input 	Instr_IF_0;
output 	Selector11;
input 	Instr_IF_1;
output 	WideOr4;
output 	WideOr41;
input 	Instr_IF_31;
output 	input_hazard_Reg_ID;
output 	WideOr21;
output 	Selector141;
output 	WideOr211;
output 	WideOr212;
output 	WideOr14;
output 	WideOr6;
output 	WideOr61;
output 	WideOr33;
output 	Decoder0;
output 	WideOr11;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Decoder0~0_combout ;
wire \Selector14~1_combout ;
wire \WideOr21~1_combout ;


// Location: LCCOMB_X56_Y28_N30
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// Selector14 = (!Instr_IF_28 & (!Instr_IF_26 & (!Instr_IF_30 & !Instr_IF_27)))

	.dataa(Instr_IF_28),
	.datab(Instr_IF_26),
	.datac(Instr_IF_30),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'h0001;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N2
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// Selector11 = (Instr_IF_29) # (!Selector14)

	.dataa(Selector14),
	.datab(gnd),
	.datac(Instr_IF_29),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hF5F5;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N10
cycloneive_lcell_comb \WideOr4~0 (
// Equation(s):
// WideOr4 = (Instr_IF_2 & ((Instr_IF_1) # ((!Instr_IF_5)))) # (!Instr_IF_2 & (((Instr_IF_0) # (Instr_IF_5))))

	.dataa(Instr_IF_1),
	.datab(Instr_IF_2),
	.datac(Instr_IF_0),
	.datad(Instr_IF_5),
	.cin(gnd),
	.combout(WideOr4),
	.cout());
// synopsys translate_off
defparam \WideOr4~0 .lut_mask = 16'hBBFC;
defparam \WideOr4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N28
cycloneive_lcell_comb \WideOr4~1 (
// Equation(s):
// WideOr41 = (!Instr_IF_1 & (!Instr_IF_2 & (!Instr_IF_0 & !Instr_IF_5)))

	.dataa(Instr_IF_1),
	.datab(Instr_IF_2),
	.datac(Instr_IF_0),
	.datad(Instr_IF_5),
	.cin(gnd),
	.combout(WideOr41),
	.cout());
// synopsys translate_off
defparam \WideOr4~1 .lut_mask = 16'h0001;
defparam \WideOr4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N12
cycloneive_lcell_comb \input_hazard_Reg_ID~0 (
// Equation(s):
// input_hazard_Reg_ID = (Instr_IF_29 & (((!Instr_IF_27) # (!Instr_IF_31)) # (!Instr_IF_26))) # (!Instr_IF_29 & ((Instr_IF_26) # ((Instr_IF_31) # (Instr_IF_27))))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_26),
	.datac(Instr_IF_31),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(input_hazard_Reg_ID),
	.cout());
// synopsys translate_off
defparam \input_hazard_Reg_ID~0 .lut_mask = 16'h7FFE;
defparam \input_hazard_Reg_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N10
cycloneive_lcell_comb \WideOr21~0 (
// Equation(s):
// WideOr21 = (Instr_IF_26 & (!Instr_IF_28 & Instr_IF_27))

	.dataa(gnd),
	.datab(Instr_IF_26),
	.datac(Instr_IF_28),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(WideOr21),
	.cout());
// synopsys translate_off
defparam \WideOr21~0 .lut_mask = 16'h0C00;
defparam \WideOr21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N10
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// Selector141 = (\Decoder0~0_combout  & (\Selector14~1_combout  & Selector14))

	.dataa(\Decoder0~0_combout ),
	.datab(\Selector14~1_combout ),
	.datac(Selector14),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector141),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'h8080;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N14
cycloneive_lcell_comb \WideOr21~2 (
// Equation(s):
// WideOr211 = (Instr_IF_29 & (!\WideOr21~1_combout )) # (!Instr_IF_29 & (((Instr_IF_31 & WideOr21))))

	.dataa(Instr_IF_29),
	.datab(\WideOr21~1_combout ),
	.datac(Instr_IF_31),
	.datad(WideOr21),
	.cin(gnd),
	.combout(WideOr211),
	.cout());
// synopsys translate_off
defparam \WideOr21~2 .lut_mask = 16'h7222;
defparam \WideOr21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \WideOr21~3 (
// Equation(s):
// WideOr212 = (WideOr211 & !Instr_IF_30)

	.dataa(gnd),
	.datab(WideOr211),
	.datac(gnd),
	.datad(Instr_IF_30),
	.cin(gnd),
	.combout(WideOr212),
	.cout());
// synopsys translate_off
defparam \WideOr21~3 .lut_mask = 16'h00CC;
defparam \WideOr21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N14
cycloneive_lcell_comb \WideOr14~0 (
// Equation(s):
// WideOr14 = (!Instr_IF_30 & (Instr_IF_29 & (!Instr_IF_31 & Instr_IF_28)))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_29),
	.datac(Instr_IF_31),
	.datad(Instr_IF_28),
	.cin(gnd),
	.combout(WideOr14),
	.cout());
// synopsys translate_off
defparam \WideOr14~0 .lut_mask = 16'h0400;
defparam \WideOr14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N12
cycloneive_lcell_comb \WideOr6~0 (
// Equation(s):
// WideOr6 = (Instr_IF_5 & (Instr_IF_3 $ (((Instr_IF_1 & !Instr_IF_2))))) # (!Instr_IF_5 & ((Instr_IF_1) # ((Instr_IF_2))))

	.dataa(Instr_IF_1),
	.datab(Instr_IF_5),
	.datac(Instr_IF_3),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(WideOr6),
	.cout());
// synopsys translate_off
defparam \WideOr6~0 .lut_mask = 16'hF36A;
defparam \WideOr6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N30
cycloneive_lcell_comb \WideOr6~1 (
// Equation(s):
// WideOr61 = (!Instr_IF_1 & (Instr_IF_5 & (!Instr_IF_3 & !Instr_IF_2)))

	.dataa(Instr_IF_1),
	.datab(Instr_IF_5),
	.datac(Instr_IF_3),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(WideOr61),
	.cout());
// synopsys translate_off
defparam \WideOr6~1 .lut_mask = 16'h0004;
defparam \WideOr6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N0
cycloneive_lcell_comb \WideOr33~0 (
// Equation(s):
// WideOr33 = (!Instr_IF_29 & ((Instr_IF_28 & (!Instr_IF_26 & !Instr_IF_27)) # (!Instr_IF_28 & ((Instr_IF_27)))))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_26),
	.datac(Instr_IF_28),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(WideOr33),
	.cout());
// synopsys translate_off
defparam \WideOr33~0 .lut_mask = 16'h0510;
defparam \WideOr33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N22
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// Decoder0 = (!Instr_IF_1 & (\Decoder0~0_combout  & Instr_IF_3))

	.dataa(Instr_IF_1),
	.datab(gnd),
	.datac(\Decoder0~0_combout ),
	.datad(Instr_IF_3),
	.cin(gnd),
	.combout(Decoder0),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h5000;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N20
cycloneive_lcell_comb \WideOr11~0 (
// Equation(s):
// WideOr11 = (!Instr_IF_29 & ((Instr_IF_28 & ((Instr_IF_27))) # (!Instr_IF_28 & (Instr_IF_26 & !Instr_IF_27))))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_26),
	.datac(Instr_IF_28),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
// synopsys translate_off
defparam \WideOr11~0 .lut_mask = 16'h5004;
defparam \WideOr11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N14
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (!Instr_IF_0 & (!Instr_IF_5 & (!Instr_IF_4 & !Instr_IF_2)))

	.dataa(Instr_IF_0),
	.datab(Instr_IF_5),
	.datac(Instr_IF_4),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h0001;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N8
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (!Instr_IF_3 & (!Instr_IF_29 & !Instr_IF_31))

	.dataa(Instr_IF_3),
	.datab(gnd),
	.datac(Instr_IF_29),
	.datad(Instr_IF_31),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'h0005;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N24
cycloneive_lcell_comb \WideOr21~1 (
// Equation(s):
// \WideOr21~1_combout  = (Instr_IF_28 & (((Instr_IF_31) # (!Instr_IF_27)) # (!Instr_IF_26))) # (!Instr_IF_28 & (Instr_IF_31 & ((!Instr_IF_27) # (!Instr_IF_26))))

	.dataa(Instr_IF_28),
	.datab(Instr_IF_26),
	.datac(Instr_IF_31),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(\WideOr21~1_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr21~1 .lut_mask = 16'hB2FA;
defparam \WideOr21~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module hazard_unit (
	MemToReg_EX,
	RegDst_EX_0,
	RegDst_EX_1,
	RegDst_EX_2,
	RegWen_EX,
	RegDst_EX_3,
	RegDst_EX_4,
	Instr_ID_16,
	hazard_Reg_ID,
	Instr_ID_17,
	always0,
	Instr_ID_18,
	Equal4,
	Instr_ID_19,
	Equal41,
	Instr_ID_20,
	Equal42,
	MemToReg_MEM,
	always01,
	RegWen_MEM,
	RegDst_MEM_0,
	output_RegWen_MEM,
	RegDst_MEM_1,
	RegDst_MEM_4,
	output_RegWen_MEM1,
	RegDst_MEM_3,
	RegDst_MEM_2,
	src2_hazard_t,
	Instr_ID_21,
	Instr_ID_22,
	always02,
	Instr_ID_24,
	Equal0,
	Instr_ID_25,
	Equal01,
	Instr_ID_23,
	always03,
	src1_hazard_t,
	src2_hazard_t1,
	src2_hazard_t2,
	devpor,
	devclrn,
	devoe);
input 	MemToReg_EX;
input 	RegDst_EX_0;
input 	RegDst_EX_1;
input 	RegDst_EX_2;
input 	RegWen_EX;
input 	RegDst_EX_3;
input 	RegDst_EX_4;
input 	Instr_ID_16;
input 	hazard_Reg_ID;
input 	Instr_ID_17;
output 	always0;
input 	Instr_ID_18;
output 	Equal4;
input 	Instr_ID_19;
output 	Equal41;
input 	Instr_ID_20;
output 	Equal42;
input 	MemToReg_MEM;
output 	always01;
input 	RegWen_MEM;
input 	RegDst_MEM_0;
input 	output_RegWen_MEM;
input 	RegDst_MEM_1;
input 	RegDst_MEM_4;
input 	output_RegWen_MEM1;
input 	RegDst_MEM_3;
input 	RegDst_MEM_2;
output 	src2_hazard_t;
input 	Instr_ID_21;
input 	Instr_ID_22;
output 	always02;
input 	Instr_ID_24;
output 	Equal0;
input 	Instr_ID_25;
output 	Equal01;
input 	Instr_ID_23;
output 	always03;
output 	src1_hazard_t;
output 	src2_hazard_t1;
output 	src2_hazard_t2;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \Equal1~1_combout ;
wire \Equal1~0_combout ;
wire \Equal5~0_combout ;
wire \src2_hazard_t~0_combout ;
wire \Equal5~2_combout ;
wire \Equal3~0_combout ;
wire \Equal3~1_combout ;
wire \Equal5~1_combout ;
wire \src2_hazard_t~1_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \always0~3_combout ;
wire \always0~4_combout ;
wire \always0~6_combout ;
wire \always0~5_combout ;
wire \always0~7_combout ;
wire \Equal2~2_combout ;
wire \Equal2~3_combout ;
wire \Equal2~1_combout ;
wire \Equal2~0_combout ;
wire \src1_hazard_t~0_combout ;


// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// always0 = (!\Equal4~0_combout  & (!\Equal4~1_combout  & ((!\Equal1~0_combout ) # (!\Equal1~1_combout ))))

	.dataa(\Equal4~0_combout ),
	.datab(\Equal4~1_combout ),
	.datac(\Equal1~1_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h0111;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Equal4~2 (
// Equation(s):
// Equal4 = (RegWen_EX1 & (RegDst_EX_2 $ (((Instr_ID_18 & hazard_Reg_ID1))))) # (!RegWen_EX1 & (Instr_ID_18 & ((hazard_Reg_ID1))))

	.dataa(RegWen_EX),
	.datab(Instr_ID_18),
	.datac(RegDst_EX_2),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(Equal4),
	.cout());
// synopsys translate_off
defparam \Equal4~2 .lut_mask = 16'h6CA0;
defparam \Equal4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Equal4~3 (
// Equation(s):
// Equal41 = (RegDst_EX_3 & (RegWen_EX1 $ (((hazard_Reg_ID1 & Instr_ID_19))))) # (!RegDst_EX_3 & (hazard_Reg_ID1 & (Instr_ID_19)))

	.dataa(RegDst_EX_3),
	.datab(hazard_Reg_ID),
	.datac(Instr_ID_19),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(Equal41),
	.cout());
// synopsys translate_off
defparam \Equal4~3 .lut_mask = 16'h6AC0;
defparam \Equal4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \Equal4~4 (
// Equation(s):
// Equal42 = (RegWen_EX1 & (RegDst_EX_4 $ (((Instr_ID_20 & hazard_Reg_ID1))))) # (!RegWen_EX1 & (((Instr_ID_20 & hazard_Reg_ID1))))

	.dataa(RegWen_EX),
	.datab(RegDst_EX_4),
	.datac(Instr_ID_20),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(Equal42),
	.cout());
// synopsys translate_off
defparam \Equal4~4 .lut_mask = 16'h7888;
defparam \Equal4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// always01 = (!Equal41 & (!Equal42 & (!Equal4 & always0)))

	.dataa(Equal41),
	.datab(Equal42),
	.datac(Equal4),
	.datad(always0),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h0100;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \src2_hazard_t~2 (
// Equation(s):
// src2_hazard_t = (\src2_hazard_t~0_combout  & (!\Equal5~2_combout  & (!\Equal3~1_combout  & \src2_hazard_t~1_combout )))

	.dataa(\src2_hazard_t~0_combout ),
	.datab(\Equal5~2_combout ),
	.datac(\Equal3~1_combout ),
	.datad(\src2_hazard_t~1_combout ),
	.cin(gnd),
	.combout(src2_hazard_t),
	.cout());
// synopsys translate_off
defparam \src2_hazard_t~2 .lut_mask = 16'h0200;
defparam \src2_hazard_t~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// always02 = (!\Equal0~0_combout  & (!\Equal0~1_combout  & ((!\Equal1~0_combout ) # (!\Equal1~1_combout ))))

	.dataa(\Equal0~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h0105;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// Equal0 = Instr_ID_24 $ (((RegDst_EX_3 & RegWen_EX1)))

	.dataa(gnd),
	.datab(Instr_ID_24),
	.datac(RegDst_EX_3),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h3CCC;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// Equal01 = Instr_ID_25 $ (((RegDst_EX_4 & RegWen_EX1)))

	.dataa(Instr_ID_25),
	.datab(RegDst_EX_4),
	.datac(gnd),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(Equal01),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'h66AA;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// always03 = (\always0~3_combout  & (\always0~7_combout  & ((!\Equal1~0_combout ) # (!\Equal1~1_combout ))))

	.dataa(\Equal1~1_combout ),
	.datab(\always0~3_combout ),
	.datac(\Equal1~0_combout ),
	.datad(\always0~7_combout ),
	.cin(gnd),
	.combout(always03),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h4C00;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \src1_hazard_t~1 (
// Equation(s):
// src1_hazard_t = (!\Equal2~2_combout  & (!\Equal2~3_combout  & (!\Equal3~1_combout  & \src1_hazard_t~0_combout )))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~3_combout ),
	.datac(\Equal3~1_combout ),
	.datad(\src1_hazard_t~0_combout ),
	.cin(gnd),
	.combout(src1_hazard_t),
	.cout());
// synopsys translate_off
defparam \src1_hazard_t~1 .lut_mask = 16'h0100;
defparam \src1_hazard_t~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \src2_hazard_t~3 (
// Equation(s):
// src2_hazard_t1 = (always01 & (((MemToReg_EX1)))) # (!always01 & (src2_hazard_t & ((!MemToReg_EX1) # (!MemToReg_MEM1))))

	.dataa(MemToReg_MEM),
	.datab(src2_hazard_t),
	.datac(always01),
	.datad(MemToReg_EX),
	.cin(gnd),
	.combout(src2_hazard_t1),
	.cout());
// synopsys translate_off
defparam \src2_hazard_t~3 .lut_mask = 16'hF40C;
defparam \src2_hazard_t~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \src2_hazard_t~4 (
// Equation(s):
// src2_hazard_t2 = (src2_hazard_t & (!always01 & (MemToReg_MEM1 & MemToReg_EX1)))

	.dataa(src2_hazard_t),
	.datab(always01),
	.datac(MemToReg_MEM),
	.datad(MemToReg_EX),
	.cin(gnd),
	.combout(src2_hazard_t2),
	.cout());
// synopsys translate_off
defparam \src2_hazard_t~4 .lut_mask = 16'h2000;
defparam \src2_hazard_t~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Equal4~0 (
// Equation(s):
// \Equal4~0_combout  = (RegWen_EX1 & (RegDst_EX_0 $ (((Instr_ID_16 & hazard_Reg_ID1))))) # (!RegWen_EX1 & (Instr_ID_16 & ((hazard_Reg_ID1))))

	.dataa(RegWen_EX),
	.datab(Instr_ID_16),
	.datac(RegDst_EX_0),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~0 .lut_mask = 16'h6CA0;
defparam \Equal4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \Equal4~1 (
// Equation(s):
// \Equal4~1_combout  = (Instr_ID_17 & (hazard_Reg_ID1 $ (((RegDst_EX_1 & RegWen_EX1))))) # (!Instr_ID_17 & (RegDst_EX_1 & (RegWen_EX1)))

	.dataa(Instr_ID_17),
	.datab(RegDst_EX_1),
	.datac(RegWen_EX),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~1 .lut_mask = 16'h6AC0;
defparam \Equal4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Equal1~1 (
// Equation(s):
// \Equal1~1_combout  = ((!RegDst_EX_4 & !RegDst_EX_3)) # (!RegWen_EX1)

	.dataa(RegDst_EX_4),
	.datab(gnd),
	.datac(RegDst_EX_3),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'h05FF;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// \Equal1~0_combout  = ((!RegDst_EX_2 & (!RegDst_EX_1 & !RegDst_EX_0))) # (!RegWen_EX1)

	.dataa(RegDst_EX_2),
	.datab(RegDst_EX_1),
	.datac(RegDst_EX_0),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h01FF;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \Equal5~0 (
// Equation(s):
// \Equal5~0_combout  = (RegWen_MEM1 & (RegDst_MEM_1 $ (((hazard_Reg_ID1 & Instr_ID_17))))) # (!RegWen_MEM1 & (hazard_Reg_ID1 & ((Instr_ID_17))))

	.dataa(RegWen_MEM),
	.datab(hazard_Reg_ID),
	.datac(RegDst_MEM_1),
	.datad(Instr_ID_17),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~0 .lut_mask = 16'h6CA0;
defparam \Equal5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \src2_hazard_t~0 (
// Equation(s):
// \src2_hazard_t~0_combout  = (!\Equal5~0_combout  & (\output_RegWen_MEM~0_combout  $ (((!Instr_ID_16) # (!hazard_Reg_ID1)))))

	.dataa(\Equal5~0_combout ),
	.datab(hazard_Reg_ID),
	.datac(output_RegWen_MEM),
	.datad(Instr_ID_16),
	.cin(gnd),
	.combout(\src2_hazard_t~0_combout ),
	.cout());
// synopsys translate_off
defparam \src2_hazard_t~0 .lut_mask = 16'h4105;
defparam \src2_hazard_t~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Equal5~2 (
// Equation(s):
// \Equal5~2_combout  = (Instr_ID_18 & (hazard_Reg_ID1 $ (((RegDst_MEM_2 & RegWen_MEM1))))) # (!Instr_ID_18 & (RegDst_MEM_2 & (RegWen_MEM1)))

	.dataa(Instr_ID_18),
	.datab(RegDst_MEM_2),
	.datac(RegWen_MEM),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(\Equal5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~2 .lut_mask = 16'h6AC0;
defparam \Equal5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = (!RegDst_MEM_3 & (!RegDst_MEM_2 & !RegDst_MEM_0))

	.dataa(gnd),
	.datab(RegDst_MEM_3),
	.datac(RegDst_MEM_2),
	.datad(RegDst_MEM_0),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0003;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// \Equal3~1_combout  = ((!RegDst_MEM_4 & (!RegDst_MEM_1 & \Equal3~0_combout ))) # (!RegWen_MEM1)

	.dataa(RegDst_MEM_4),
	.datab(RegDst_MEM_1),
	.datac(RegWen_MEM),
	.datad(\Equal3~0_combout ),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h1F0F;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Equal5~1 (
// Equation(s):
// \Equal5~1_combout  = (RegWen_MEM1 & (RegDst_MEM_3 $ (((Instr_ID_19 & hazard_Reg_ID1))))) # (!RegWen_MEM1 & (Instr_ID_19 & ((hazard_Reg_ID1))))

	.dataa(RegWen_MEM),
	.datab(Instr_ID_19),
	.datac(RegDst_MEM_3),
	.datad(hazard_Reg_ID),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~1 .lut_mask = 16'h6CA0;
defparam \Equal5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \src2_hazard_t~1 (
// Equation(s):
// \src2_hazard_t~1_combout  = (!\Equal5~1_combout  & (\output_RegWen_MEM~1_combout  $ (((!Instr_ID_20) # (!hazard_Reg_ID1)))))

	.dataa(\Equal5~1_combout ),
	.datab(hazard_Reg_ID),
	.datac(Instr_ID_20),
	.datad(output_RegWen_MEM1),
	.cin(gnd),
	.combout(\src2_hazard_t~1_combout ),
	.cout());
// synopsys translate_off
defparam \src2_hazard_t~1 .lut_mask = 16'h4015;
defparam \src2_hazard_t~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = Instr_ID_21 $ (((RegDst_EX_0 & RegWen_EX1)))

	.dataa(RegDst_EX_0),
	.datab(Instr_ID_21),
	.datac(gnd),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h66CC;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = Instr_ID_22 $ (((RegDst_EX_1 & RegWen_EX1)))

	.dataa(gnd),
	.datab(RegDst_EX_1),
	.datac(Instr_ID_22),
	.datad(RegWen_EX),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h3CF0;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (RegWen_EX1 & (Instr_ID_24 $ ((!RegDst_EX_3)))) # (!RegWen_EX1 & (!Instr_ID_24 & ((!Instr_ID_21))))

	.dataa(Instr_ID_24),
	.datab(RegWen_EX),
	.datac(RegDst_EX_3),
	.datad(Instr_ID_21),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h8495;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (RegDst_EX_0 & (Instr_ID_21 & (RegDst_EX_1 $ (!Instr_ID_22)))) # (!RegDst_EX_0 & (!Instr_ID_21 & (RegDst_EX_1 $ (!Instr_ID_22))))

	.dataa(RegDst_EX_0),
	.datab(RegDst_EX_1),
	.datac(Instr_ID_21),
	.datad(Instr_ID_22),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8421;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (!Instr_ID_25 & (!Instr_ID_23 & !Instr_ID_22))

	.dataa(gnd),
	.datab(Instr_ID_25),
	.datac(Instr_ID_23),
	.datad(Instr_ID_22),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'h0003;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (RegDst_EX_2 & (Instr_ID_23 & (Instr_ID_25 $ (!RegDst_EX_4)))) # (!RegDst_EX_2 & (!Instr_ID_23 & (Instr_ID_25 $ (!RegDst_EX_4))))

	.dataa(RegDst_EX_2),
	.datab(Instr_ID_25),
	.datac(Instr_ID_23),
	.datad(RegDst_EX_4),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8421;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (RegWen_EX1 & (\always0~4_combout  & ((\always0~5_combout )))) # (!RegWen_EX1 & (((\always0~6_combout ))))

	.dataa(RegWen_EX),
	.datab(\always0~4_combout ),
	.datac(\always0~6_combout ),
	.datad(\always0~5_combout ),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'hD850;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = Instr_ID_21 $ (((RegDst_MEM_0 & RegWen_MEM1)))

	.dataa(gnd),
	.datab(RegDst_MEM_0),
	.datac(Instr_ID_21),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h3CF0;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = Instr_ID_22 $ (((RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(gnd),
	.datab(Instr_ID_22),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h3CCC;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = Instr_ID_24 $ (((RegWen_MEM1 & RegDst_MEM_3)))

	.dataa(RegWen_MEM),
	.datab(RegDst_MEM_3),
	.datac(gnd),
	.datad(Instr_ID_24),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h7788;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = Instr_ID_23 $ (((RegWen_MEM1 & RegDst_MEM_2)))

	.dataa(gnd),
	.datab(RegWen_MEM),
	.datac(Instr_ID_23),
	.datad(RegDst_MEM_2),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h3CF0;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \src1_hazard_t~0 (
// Equation(s):
// \src1_hazard_t~0_combout  = (!\Equal2~1_combout  & (!\Equal2~0_combout  & (\output_RegWen_MEM~1_combout  $ (!Instr_ID_25))))

	.dataa(output_RegWen_MEM1),
	.datab(Instr_ID_25),
	.datac(\Equal2~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\src1_hazard_t~0_combout ),
	.cout());
// synopsys translate_off
defparam \src1_hazard_t~0 .lut_mask = 16'h0009;
defparam \src1_hazard_t~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_registers (
	pc_next_plus4_2,
	pc_next_plus4_3,
	pc_next_plus4_4,
	pc_next_plus4_5,
	pc_next_plus4_6,
	pc_next_plus4_7,
	pc_next_plus4_8,
	pc_next_plus4_9,
	pc_next_plus4_10,
	pc_next_plus4_11,
	pc_next_plus4_12,
	pc_next_plus4_13,
	pc_next_plus4_14,
	pc_next_plus4_15,
	pc_next_plus4_16,
	pc_next_plus4_17,
	pc_next_plus4_18,
	pc_next_plus4_19,
	pc_next_plus4_20,
	pc_next_plus4_21,
	pc_next_plus4_22,
	pc_next_plus4_23,
	pc_next_plus4_24,
	pc_next_plus4_25,
	pc_next_plus4_26,
	pc_next_plus4_27,
	pc_next_plus4_28,
	pc_next_plus4_29,
	pc_next_plus4_30,
	pc_next_plus4_31,
	Result_EX_1,
	pc_1,
	Memwrite_EX1,
	MemToReg_EX1,
	Result_EX_0,
	pc_0,
	Result_EX_3,
	Result_EX_2,
	Result_EX_5,
	Result_EX_4,
	Result_EX_7,
	Result_EX_6,
	Result_EX_9,
	Result_EX_8,
	Result_EX_11,
	Result_EX_10,
	Result_EX_13,
	Result_EX_12,
	Result_EX_15,
	Result_EX_14,
	Result_EX_17,
	Result_EX_16,
	Result_EX_19,
	Result_EX_18,
	Result_EX_21,
	Result_EX_20,
	Result_EX_23,
	Result_EX_22,
	Result_EX_25,
	Result_EX_24,
	Result_EX_27,
	Result_EX_26,
	Result_EX_29,
	Result_EX_28,
	Result_EX_31,
	Result_EX_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	halt_MEM1,
	care_ID1,
	ALUOP_ID_1,
	ALUOP_ID_3,
	ALUOP_ID_2,
	RegDst_EX_0,
	RegDst_EX_1,
	RegDst_EX_2,
	RegWen_EX1,
	RegDst_EX_3,
	RegDst_EX_4,
	Instr_ID_16,
	hazard_Reg_ID1,
	Instr_ID_17,
	Instr_ID_18,
	Instr_ID_19,
	Memwrite_ID1,
	Instr_ID_20,
	ReadData_MEM_31,
	CalcData_MEM_31,
	MemToReg_MEM1,
	input_a,
	always0,
	RegWen_MEM1,
	RegDst_MEM_0,
	RegDst_MEM_1,
	RegDst_MEM_4,
	RegDst_MEM_3,
	RegDst_MEM_2,
	ALUSrc2_ID_31,
	Instr_ID_21,
	Instr_ID_22,
	Instr_ID_24,
	Instr_ID_25,
	Instr_ID_23,
	ALUSrc1_ID_31,
	always01,
	src1_hazard_t,
	ALUOP_ID_0,
	ALUSrc1_ID_30,
	ReadData_MEM_30,
	CalcData_MEM_30,
	input_b,
	ALUSrc2_ID_30,
	ALUSrc1_ID_29,
	ReadData_MEM_29,
	CalcData_MEM_29,
	input_b1,
	ALUSrc2_ID_29,
	ALUSrc1_ID_28,
	ReadData_MEM_28,
	CalcData_MEM_28,
	input_b2,
	ALUSrc2_ID_28,
	ALUSrc1_ID_27,
	ReadData_MEM_27,
	CalcData_MEM_27,
	input_b3,
	ALUSrc2_ID_27,
	ALUSrc1_ID_26,
	ReadData_MEM_26,
	CalcData_MEM_26,
	input_b4,
	ALUSrc2_ID_26,
	ALUSrc1_ID_25,
	ReadData_MEM_25,
	CalcData_MEM_25,
	input_b5,
	ALUSrc2_ID_25,
	ALUSrc1_ID_24,
	ReadData_MEM_24,
	CalcData_MEM_24,
	input_b6,
	ALUSrc2_ID_24,
	ALUSrc1_ID_23,
	ReadData_MEM_23,
	CalcData_MEM_23,
	input_b7,
	ALUSrc2_ID_23,
	ALUSrc1_ID_22,
	ReadData_MEM_22,
	CalcData_MEM_22,
	input_b8,
	ALUSrc2_ID_22,
	ALUSrc1_ID_21,
	ReadData_MEM_21,
	CalcData_MEM_21,
	input_b9,
	ALUSrc2_ID_21,
	ALUSrc1_ID_20,
	ReadData_MEM_20,
	CalcData_MEM_20,
	input_b10,
	ALUSrc2_ID_20,
	ALUSrc1_ID_19,
	ReadData_MEM_19,
	CalcData_MEM_19,
	input_b11,
	ALUSrc2_ID_19,
	ALUSrc1_ID_18,
	ReadData_MEM_18,
	CalcData_MEM_18,
	input_b12,
	ALUSrc2_ID_18,
	ALUSrc1_ID_17,
	ReadData_MEM_17,
	CalcData_MEM_17,
	input_b13,
	ALUSrc2_ID_17,
	ALUSrc1_ID_16,
	ReadData_MEM_16,
	CalcData_MEM_16,
	input_b14,
	ALUSrc2_ID_16,
	ALUSrc1_ID_15,
	ReadData_MEM_15,
	CalcData_MEM_15,
	input_b15,
	ALUSrc2_ID_15,
	ALUSrc1_ID_14,
	ReadData_MEM_14,
	CalcData_MEM_14,
	input_b16,
	ALUSrc2_ID_14,
	ReadData_MEM_13,
	CalcData_MEM_13,
	input_a1,
	ALUSrc2_ID_13,
	ALUSrc1_ID_13,
	ReadData_MEM_12,
	CalcData_MEM_12,
	input_a2,
	ALUSrc2_ID_12,
	ALUSrc1_ID_12,
	ReadData_MEM_11,
	CalcData_MEM_11,
	input_a3,
	ALUSrc2_ID_11,
	ALUSrc1_ID_11,
	ReadData_MEM_10,
	CalcData_MEM_10,
	input_a4,
	ALUSrc2_ID_10,
	ALUSrc1_ID_10,
	ReadData_MEM_9,
	CalcData_MEM_9,
	input_a5,
	ALUSrc2_ID_9,
	ALUSrc1_ID_9,
	ReadData_MEM_8,
	CalcData_MEM_8,
	input_a6,
	ALUSrc2_ID_8,
	ALUSrc1_ID_8,
	ReadData_MEM_7,
	CalcData_MEM_7,
	input_a7,
	ALUSrc2_ID_7,
	ALUSrc1_ID_7,
	ReadData_MEM_6,
	CalcData_MEM_6,
	input_a8,
	ALUSrc2_ID_6,
	ALUSrc1_ID_6,
	ReadData_MEM_5,
	CalcData_MEM_5,
	input_a9,
	ALUSrc2_ID_5,
	ALUSrc1_ID_5,
	ReadData_MEM_4,
	CalcData_MEM_4,
	input_a10,
	ALUSrc2_ID_4,
	ALUSrc1_ID_4,
	ReadData_MEM_3,
	CalcData_MEM_3,
	input_a11,
	ALUSrc2_ID_3,
	ALUSrc1_ID_3,
	ReadData_MEM_2,
	CalcData_MEM_2,
	input_a12,
	ALUSrc2_ID_2,
	ALUSrc1_ID_2,
	ReadData_MEM_1,
	CalcData_MEM_1,
	input_a13,
	ALUSrc2_ID_1,
	ALUSrc1_ID_1,
	ReadData_MEM_0,
	CalcData_MEM_0,
	input_a14,
	ALUSrc2_ID_0,
	ALUSrc1_ID_0,
	Wdata_EX_0,
	src2_hazard_t,
	nextPC_ID_1,
	Selector30,
	jump_ID_0,
	jump_ID_1,
	jump_ID_2,
	Equal8,
	Selector28,
	Selector3,
	Selector22,
	Selector2,
	Selector27,
	Selector25,
	Selector24,
	Selector26,
	Selector4,
	Selector16,
	Selector7,
	Selector6,
	Selector29,
	Selector15,
	Selector5,
	Selector31,
	Selector11,
	Selector10,
	Selector21,
	Selector20,
	Selector9,
	Selector8,
	Selector14,
	Selector13,
	Selector12,
	Selector23,
	Selector19,
	Selector18,
	Selector17,
	Selector0,
	Selector1,
	branch,
	always02,
	nextPC_ID_0,
	nextPC_ID_3,
	Instr_ID_1,
	nextPC_ID_2,
	Instr_ID_0,
	nextPC_ID_5,
	Instr_ID_3,
	nextPC_ID_4,
	Instr_ID_2,
	nextPC_ID_7,
	Instr_ID_5,
	nextPC_ID_6,
	Instr_ID_4,
	nextPC_ID_9,
	Instr_ID_7,
	nextPC_ID_8,
	Instr_ID_6,
	nextPC_ID_11,
	Instr_ID_9,
	nextPC_ID_10,
	Instr_ID_8,
	nextPC_ID_13,
	Instr_ID_11,
	nextPC_ID_12,
	Instr_ID_10,
	nextPC_ID_15,
	Instr_ID_13,
	nextPC_ID_14,
	Instr_ID_12,
	nextPC_ID_17,
	Instr_ID_15,
	nextPC_ID_16,
	Instr_ID_14,
	nextPC_ID_19,
	nextPC_ID_18,
	nextPC_ID_21,
	nextPC_ID_20,
	nextPC_ID_23,
	nextPC_ID_22,
	nextPC_ID_25,
	nextPC_ID_24,
	nextPC_ID_27,
	nextPC_ID_26,
	nextPC_ID_29,
	nextPC_ID_28,
	nextPC_ID_31,
	nextPC_ID_30,
	Wdata_EX_1,
	Wdata_EX_2,
	Wdata_EX_3,
	Wdata_EX_4,
	Wdata_EX_5,
	Wdata_EX_6,
	Wdata_EX_7,
	Wdata_EX_8,
	Wdata_EX_9,
	Wdata_EX_10,
	Wdata_EX_11,
	Wdata_EX_12,
	Wdata_EX_13,
	Wdata_EX_14,
	Wdata_EX_15,
	Wdata_EX_16,
	Wdata_EX_17,
	Wdata_EX_18,
	Wdata_EX_19,
	Wdata_EX_20,
	Wdata_EX_21,
	Wdata_EX_22,
	Wdata_EX_23,
	Wdata_EX_24,
	Wdata_EX_25,
	Wdata_EX_26,
	Wdata_EX_27,
	Wdata_EX_28,
	Wdata_EX_29,
	Wdata_EX_30,
	Wdata_EX_31,
	Instr_IF_30,
	Instr_IF_28,
	Instr_IF_26,
	Instr_IF_27,
	Selector141,
	Instr_IF_29,
	Instr_IF_5,
	Instr_IF_4,
	Instr_IF_2,
	Instr_IF_3,
	Instr_IF_0,
	src2_hazard_t1,
	Selector111,
	Instr_IF_1,
	WideOr4,
	WideOr41,
	Instr_IF_31,
	Instr_IF_16,
	input_hazard_Reg_ID,
	Instr_IF_17,
	Instr_IF_18,
	Instr_IF_19,
	WideOr21,
	Instr_IF_20,
	Equal20,
	Selector142,
	WideOr211,
	WideOr212,
	rfifrdat2_31,
	WideOr14,
	Instr_IF_21,
	Instr_IF_22,
	Instr_IF_24,
	Instr_IF_25,
	Instr_IF_23,
	rfifrdat1_31,
	rfifrdat1_311,
	WideOr0,
	WideOr6,
	WideOr61,
	rfifrdat1_30,
	rfifrdat1_301,
	rfifrdat2_30,
	rfifrdat1_29,
	rfifrdat1_291,
	rfifrdat2_29,
	rfifrdat1_28,
	rfifrdat1_281,
	rfifrdat2_28,
	rfifrdat1_27,
	rfifrdat1_271,
	rfifrdat2_27,
	rfifrdat1_26,
	rfifrdat1_261,
	rfifrdat2_26,
	Instr_IF_10,
	rfifrdat1_25,
	rfifrdat1_251,
	rfifrdat2_25,
	Instr_IF_9,
	rfifrdat1_24,
	rfifrdat1_241,
	rfifrdat2_24,
	Instr_IF_8,
	rfifrdat1_23,
	rfifrdat1_231,
	rfifrdat2_23,
	Instr_IF_7,
	rfifrdat1_22,
	rfifrdat1_221,
	rfifrdat2_22,
	Instr_IF_6,
	rfifrdat1_21,
	rfifrdat1_211,
	rfifrdat2_21,
	rfifrdat1_20,
	rfifrdat1_201,
	rfifrdat2_20,
	rfifrdat1_19,
	rfifrdat1_191,
	rfifrdat2_19,
	rfifrdat1_18,
	rfifrdat1_181,
	rfifrdat2_18,
	rfifrdat1_17,
	rfifrdat1_171,
	rfifrdat2_17,
	rfifrdat1_16,
	rfifrdat1_161,
	rfifrdat2_16,
	rfifrdat1_15,
	rfifrdat1_151,
	Equal0,
	rfifrdat2_15,
	rfifrdat1_14,
	rfifrdat1_141,
	rfifrdat2_14,
	rfifrdat2_13,
	rfifrdat1_13,
	rfifrdat1_131,
	rfifrdat2_12,
	rfifrdat1_12,
	rfifrdat1_121,
	rfifrdat2_11,
	rfifrdat1_11,
	rfifrdat1_111,
	rfifrdat2_10,
	rfifrdat1_10,
	rfifrdat1_101,
	rfifrdat2_9,
	rfifrdat1_9,
	rfifrdat1_91,
	rfifrdat2_8,
	rfifrdat1_8,
	rfifrdat1_81,
	rfifrdat2_7,
	rfifrdat1_7,
	rfifrdat1_71,
	rfifrdat2_6,
	rfifrdat1_6,
	rfifrdat1_61,
	rfifrdat2_5,
	rfifrdat1_5,
	rfifrdat1_51,
	rfifrdat2_4,
	input_ALUSrc2_ID,
	rfifrdat1_4,
	rfifrdat1_41,
	rfifrdat2_3,
	input_ALUSrc2_ID1,
	rfifrdat1_3,
	rfifrdat1_32,
	rfifrdat2_2,
	input_ALUSrc2_ID2,
	rfifrdat1_2,
	rfifrdat1_210,
	rfifrdat2_1,
	input_ALUSrc2_ID3,
	rfifrdat1_1,
	rfifrdat1_110,
	rfifrdat2_0,
	input_ALUSrc2_ID4,
	rfifrdat1_0,
	rfifrdat1_01,
	Equal27,
	WideOr33,
	Decoder0,
	WideOr11,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	pc_next_plus4_2;
input 	pc_next_plus4_3;
input 	pc_next_plus4_4;
input 	pc_next_plus4_5;
input 	pc_next_plus4_6;
input 	pc_next_plus4_7;
input 	pc_next_plus4_8;
input 	pc_next_plus4_9;
input 	pc_next_plus4_10;
input 	pc_next_plus4_11;
input 	pc_next_plus4_12;
input 	pc_next_plus4_13;
input 	pc_next_plus4_14;
input 	pc_next_plus4_15;
input 	pc_next_plus4_16;
input 	pc_next_plus4_17;
input 	pc_next_plus4_18;
input 	pc_next_plus4_19;
input 	pc_next_plus4_20;
input 	pc_next_plus4_21;
input 	pc_next_plus4_22;
input 	pc_next_plus4_23;
input 	pc_next_plus4_24;
input 	pc_next_plus4_25;
input 	pc_next_plus4_26;
input 	pc_next_plus4_27;
input 	pc_next_plus4_28;
input 	pc_next_plus4_29;
input 	pc_next_plus4_30;
input 	pc_next_plus4_31;
output 	Result_EX_1;
input 	pc_1;
output 	Memwrite_EX1;
output 	MemToReg_EX1;
output 	Result_EX_0;
input 	pc_0;
output 	Result_EX_3;
output 	Result_EX_2;
output 	Result_EX_5;
output 	Result_EX_4;
output 	Result_EX_7;
output 	Result_EX_6;
output 	Result_EX_9;
output 	Result_EX_8;
output 	Result_EX_11;
output 	Result_EX_10;
output 	Result_EX_13;
output 	Result_EX_12;
output 	Result_EX_15;
output 	Result_EX_14;
output 	Result_EX_17;
output 	Result_EX_16;
output 	Result_EX_19;
output 	Result_EX_18;
output 	Result_EX_21;
output 	Result_EX_20;
output 	Result_EX_23;
output 	Result_EX_22;
output 	Result_EX_25;
output 	Result_EX_24;
output 	Result_EX_27;
output 	Result_EX_26;
output 	Result_EX_29;
output 	Result_EX_28;
output 	Result_EX_31;
output 	Result_EX_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	halt_MEM1;
output 	care_ID1;
output 	ALUOP_ID_1;
output 	ALUOP_ID_3;
output 	ALUOP_ID_2;
output 	RegDst_EX_0;
output 	RegDst_EX_1;
output 	RegDst_EX_2;
output 	RegWen_EX1;
output 	RegDst_EX_3;
output 	RegDst_EX_4;
output 	Instr_ID_16;
output 	hazard_Reg_ID1;
output 	Instr_ID_17;
output 	Instr_ID_18;
output 	Instr_ID_19;
output 	Memwrite_ID1;
output 	Instr_ID_20;
output 	ReadData_MEM_31;
output 	CalcData_MEM_31;
output 	MemToReg_MEM1;
input 	input_a;
input 	always0;
output 	RegWen_MEM1;
output 	RegDst_MEM_0;
output 	RegDst_MEM_1;
output 	RegDst_MEM_4;
output 	RegDst_MEM_3;
output 	RegDst_MEM_2;
output 	ALUSrc2_ID_31;
output 	Instr_ID_21;
output 	Instr_ID_22;
output 	Instr_ID_24;
output 	Instr_ID_25;
output 	Instr_ID_23;
output 	ALUSrc1_ID_31;
input 	always01;
input 	src1_hazard_t;
output 	ALUOP_ID_0;
output 	ALUSrc1_ID_30;
output 	ReadData_MEM_30;
output 	CalcData_MEM_30;
input 	input_b;
output 	ALUSrc2_ID_30;
output 	ALUSrc1_ID_29;
output 	ReadData_MEM_29;
output 	CalcData_MEM_29;
input 	input_b1;
output 	ALUSrc2_ID_29;
output 	ALUSrc1_ID_28;
output 	ReadData_MEM_28;
output 	CalcData_MEM_28;
input 	input_b2;
output 	ALUSrc2_ID_28;
output 	ALUSrc1_ID_27;
output 	ReadData_MEM_27;
output 	CalcData_MEM_27;
input 	input_b3;
output 	ALUSrc2_ID_27;
output 	ALUSrc1_ID_26;
output 	ReadData_MEM_26;
output 	CalcData_MEM_26;
input 	input_b4;
output 	ALUSrc2_ID_26;
output 	ALUSrc1_ID_25;
output 	ReadData_MEM_25;
output 	CalcData_MEM_25;
input 	input_b5;
output 	ALUSrc2_ID_25;
output 	ALUSrc1_ID_24;
output 	ReadData_MEM_24;
output 	CalcData_MEM_24;
input 	input_b6;
output 	ALUSrc2_ID_24;
output 	ALUSrc1_ID_23;
output 	ReadData_MEM_23;
output 	CalcData_MEM_23;
input 	input_b7;
output 	ALUSrc2_ID_23;
output 	ALUSrc1_ID_22;
output 	ReadData_MEM_22;
output 	CalcData_MEM_22;
input 	input_b8;
output 	ALUSrc2_ID_22;
output 	ALUSrc1_ID_21;
output 	ReadData_MEM_21;
output 	CalcData_MEM_21;
input 	input_b9;
output 	ALUSrc2_ID_21;
output 	ALUSrc1_ID_20;
output 	ReadData_MEM_20;
output 	CalcData_MEM_20;
input 	input_b10;
output 	ALUSrc2_ID_20;
output 	ALUSrc1_ID_19;
output 	ReadData_MEM_19;
output 	CalcData_MEM_19;
input 	input_b11;
output 	ALUSrc2_ID_19;
output 	ALUSrc1_ID_18;
output 	ReadData_MEM_18;
output 	CalcData_MEM_18;
input 	input_b12;
output 	ALUSrc2_ID_18;
output 	ALUSrc1_ID_17;
output 	ReadData_MEM_17;
output 	CalcData_MEM_17;
input 	input_b13;
output 	ALUSrc2_ID_17;
output 	ALUSrc1_ID_16;
output 	ReadData_MEM_16;
output 	CalcData_MEM_16;
input 	input_b14;
output 	ALUSrc2_ID_16;
output 	ALUSrc1_ID_15;
output 	ReadData_MEM_15;
output 	CalcData_MEM_15;
input 	input_b15;
output 	ALUSrc2_ID_15;
output 	ALUSrc1_ID_14;
output 	ReadData_MEM_14;
output 	CalcData_MEM_14;
input 	input_b16;
output 	ALUSrc2_ID_14;
output 	ReadData_MEM_13;
output 	CalcData_MEM_13;
input 	input_a1;
output 	ALUSrc2_ID_13;
output 	ALUSrc1_ID_13;
output 	ReadData_MEM_12;
output 	CalcData_MEM_12;
input 	input_a2;
output 	ALUSrc2_ID_12;
output 	ALUSrc1_ID_12;
output 	ReadData_MEM_11;
output 	CalcData_MEM_11;
input 	input_a3;
output 	ALUSrc2_ID_11;
output 	ALUSrc1_ID_11;
output 	ReadData_MEM_10;
output 	CalcData_MEM_10;
input 	input_a4;
output 	ALUSrc2_ID_10;
output 	ALUSrc1_ID_10;
output 	ReadData_MEM_9;
output 	CalcData_MEM_9;
input 	input_a5;
output 	ALUSrc2_ID_9;
output 	ALUSrc1_ID_9;
output 	ReadData_MEM_8;
output 	CalcData_MEM_8;
input 	input_a6;
output 	ALUSrc2_ID_8;
output 	ALUSrc1_ID_8;
output 	ReadData_MEM_7;
output 	CalcData_MEM_7;
input 	input_a7;
output 	ALUSrc2_ID_7;
output 	ALUSrc1_ID_7;
output 	ReadData_MEM_6;
output 	CalcData_MEM_6;
input 	input_a8;
output 	ALUSrc2_ID_6;
output 	ALUSrc1_ID_6;
output 	ReadData_MEM_5;
output 	CalcData_MEM_5;
input 	input_a9;
output 	ALUSrc2_ID_5;
output 	ALUSrc1_ID_5;
output 	ReadData_MEM_4;
output 	CalcData_MEM_4;
input 	input_a10;
output 	ALUSrc2_ID_4;
output 	ALUSrc1_ID_4;
output 	ReadData_MEM_3;
output 	CalcData_MEM_3;
input 	input_a11;
output 	ALUSrc2_ID_3;
output 	ALUSrc1_ID_3;
output 	ReadData_MEM_2;
output 	CalcData_MEM_2;
input 	input_a12;
output 	ALUSrc2_ID_2;
output 	ALUSrc1_ID_2;
output 	ReadData_MEM_1;
output 	CalcData_MEM_1;
input 	input_a13;
output 	ALUSrc2_ID_1;
output 	ALUSrc1_ID_1;
output 	ReadData_MEM_0;
output 	CalcData_MEM_0;
input 	input_a14;
output 	ALUSrc2_ID_0;
output 	ALUSrc1_ID_0;
output 	Wdata_EX_0;
input 	src2_hazard_t;
output 	nextPC_ID_1;
input 	Selector30;
output 	jump_ID_0;
output 	jump_ID_1;
output 	jump_ID_2;
input 	Equal8;
input 	Selector28;
input 	Selector3;
input 	Selector22;
input 	Selector2;
input 	Selector27;
input 	Selector25;
input 	Selector24;
input 	Selector26;
input 	Selector4;
input 	Selector16;
input 	Selector7;
input 	Selector6;
input 	Selector29;
input 	Selector15;
input 	Selector5;
input 	Selector31;
input 	Selector11;
input 	Selector10;
input 	Selector21;
input 	Selector20;
input 	Selector9;
input 	Selector8;
input 	Selector14;
input 	Selector13;
input 	Selector12;
input 	Selector23;
input 	Selector19;
input 	Selector18;
input 	Selector17;
input 	Selector0;
input 	Selector1;
input 	branch;
input 	always02;
output 	nextPC_ID_0;
output 	nextPC_ID_3;
output 	Instr_ID_1;
output 	nextPC_ID_2;
output 	Instr_ID_0;
output 	nextPC_ID_5;
output 	Instr_ID_3;
output 	nextPC_ID_4;
output 	Instr_ID_2;
output 	nextPC_ID_7;
output 	Instr_ID_5;
output 	nextPC_ID_6;
output 	Instr_ID_4;
output 	nextPC_ID_9;
output 	Instr_ID_7;
output 	nextPC_ID_8;
output 	Instr_ID_6;
output 	nextPC_ID_11;
output 	Instr_ID_9;
output 	nextPC_ID_10;
output 	Instr_ID_8;
output 	nextPC_ID_13;
output 	Instr_ID_11;
output 	nextPC_ID_12;
output 	Instr_ID_10;
output 	nextPC_ID_15;
output 	Instr_ID_13;
output 	nextPC_ID_14;
output 	Instr_ID_12;
output 	nextPC_ID_17;
output 	Instr_ID_15;
output 	nextPC_ID_16;
output 	Instr_ID_14;
output 	nextPC_ID_19;
output 	nextPC_ID_18;
output 	nextPC_ID_21;
output 	nextPC_ID_20;
output 	nextPC_ID_23;
output 	nextPC_ID_22;
output 	nextPC_ID_25;
output 	nextPC_ID_24;
output 	nextPC_ID_27;
output 	nextPC_ID_26;
output 	nextPC_ID_29;
output 	nextPC_ID_28;
output 	nextPC_ID_31;
output 	nextPC_ID_30;
output 	Wdata_EX_1;
output 	Wdata_EX_2;
output 	Wdata_EX_3;
output 	Wdata_EX_4;
output 	Wdata_EX_5;
output 	Wdata_EX_6;
output 	Wdata_EX_7;
output 	Wdata_EX_8;
output 	Wdata_EX_9;
output 	Wdata_EX_10;
output 	Wdata_EX_11;
output 	Wdata_EX_12;
output 	Wdata_EX_13;
output 	Wdata_EX_14;
output 	Wdata_EX_15;
output 	Wdata_EX_16;
output 	Wdata_EX_17;
output 	Wdata_EX_18;
output 	Wdata_EX_19;
output 	Wdata_EX_20;
output 	Wdata_EX_21;
output 	Wdata_EX_22;
output 	Wdata_EX_23;
output 	Wdata_EX_24;
output 	Wdata_EX_25;
output 	Wdata_EX_26;
output 	Wdata_EX_27;
output 	Wdata_EX_28;
output 	Wdata_EX_29;
output 	Wdata_EX_30;
output 	Wdata_EX_31;
output 	Instr_IF_30;
output 	Instr_IF_28;
output 	Instr_IF_26;
output 	Instr_IF_27;
input 	Selector141;
output 	Instr_IF_29;
output 	Instr_IF_5;
output 	Instr_IF_4;
output 	Instr_IF_2;
output 	Instr_IF_3;
output 	Instr_IF_0;
input 	src2_hazard_t1;
input 	Selector111;
output 	Instr_IF_1;
input 	WideOr4;
input 	WideOr41;
output 	Instr_IF_31;
output 	Instr_IF_16;
input 	input_hazard_Reg_ID;
output 	Instr_IF_17;
output 	Instr_IF_18;
output 	Instr_IF_19;
input 	WideOr21;
output 	Instr_IF_20;
input 	Equal20;
input 	Selector142;
input 	WideOr211;
input 	WideOr212;
input 	rfifrdat2_31;
input 	WideOr14;
output 	Instr_IF_21;
output 	Instr_IF_22;
output 	Instr_IF_24;
output 	Instr_IF_25;
output 	Instr_IF_23;
input 	rfifrdat1_31;
input 	rfifrdat1_311;
input 	WideOr0;
input 	WideOr6;
input 	WideOr61;
input 	rfifrdat1_30;
input 	rfifrdat1_301;
input 	rfifrdat2_30;
input 	rfifrdat1_29;
input 	rfifrdat1_291;
input 	rfifrdat2_29;
input 	rfifrdat1_28;
input 	rfifrdat1_281;
input 	rfifrdat2_28;
input 	rfifrdat1_27;
input 	rfifrdat1_271;
input 	rfifrdat2_27;
input 	rfifrdat1_26;
input 	rfifrdat1_261;
input 	rfifrdat2_26;
output 	Instr_IF_10;
input 	rfifrdat1_25;
input 	rfifrdat1_251;
input 	rfifrdat2_25;
output 	Instr_IF_9;
input 	rfifrdat1_24;
input 	rfifrdat1_241;
input 	rfifrdat2_24;
output 	Instr_IF_8;
input 	rfifrdat1_23;
input 	rfifrdat1_231;
input 	rfifrdat2_23;
output 	Instr_IF_7;
input 	rfifrdat1_22;
input 	rfifrdat1_221;
input 	rfifrdat2_22;
output 	Instr_IF_6;
input 	rfifrdat1_21;
input 	rfifrdat1_211;
input 	rfifrdat2_21;
input 	rfifrdat1_20;
input 	rfifrdat1_201;
input 	rfifrdat2_20;
input 	rfifrdat1_19;
input 	rfifrdat1_191;
input 	rfifrdat2_19;
input 	rfifrdat1_18;
input 	rfifrdat1_181;
input 	rfifrdat2_18;
input 	rfifrdat1_17;
input 	rfifrdat1_171;
input 	rfifrdat2_17;
input 	rfifrdat1_16;
input 	rfifrdat1_161;
input 	rfifrdat2_16;
input 	rfifrdat1_15;
input 	rfifrdat1_151;
input 	Equal0;
input 	rfifrdat2_15;
input 	rfifrdat1_14;
input 	rfifrdat1_141;
input 	rfifrdat2_14;
input 	rfifrdat2_13;
input 	rfifrdat1_13;
input 	rfifrdat1_131;
input 	rfifrdat2_12;
input 	rfifrdat1_12;
input 	rfifrdat1_121;
input 	rfifrdat2_11;
input 	rfifrdat1_11;
input 	rfifrdat1_111;
input 	rfifrdat2_10;
input 	rfifrdat1_10;
input 	rfifrdat1_101;
input 	rfifrdat2_9;
input 	rfifrdat1_9;
input 	rfifrdat1_91;
input 	rfifrdat2_8;
input 	rfifrdat1_8;
input 	rfifrdat1_81;
input 	rfifrdat2_7;
input 	rfifrdat1_7;
input 	rfifrdat1_71;
input 	rfifrdat2_6;
input 	rfifrdat1_6;
input 	rfifrdat1_61;
input 	rfifrdat2_5;
input 	rfifrdat1_5;
input 	rfifrdat1_51;
input 	rfifrdat2_4;
input 	input_ALUSrc2_ID;
input 	rfifrdat1_4;
input 	rfifrdat1_41;
input 	rfifrdat2_3;
input 	input_ALUSrc2_ID1;
input 	rfifrdat1_3;
input 	rfifrdat1_32;
input 	rfifrdat2_2;
input 	input_ALUSrc2_ID2;
input 	rfifrdat1_2;
input 	rfifrdat1_210;
input 	rfifrdat2_1;
input 	input_ALUSrc2_ID3;
input 	rfifrdat1_1;
input 	rfifrdat1_110;
input 	rfifrdat2_0;
input 	input_ALUSrc2_ID4;
input 	rfifrdat1_0;
input 	rfifrdat1_01;
input 	Equal27;
input 	WideOr33;
input 	Decoder0;
input 	WideOr11;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \RegWen_ID~0_combout ;
wire \RegWen_ID~1_combout ;
wire \RegDat2_ID~0_combout ;
wire \RegDat2_ID~3_combout ;
wire \RegDat2_ID~4_combout ;
wire \RegDat2_ID~13_combout ;
wire \RegDat2_ID~17_combout ;
wire \RegDat2_ID~22_combout ;
wire \RegDat2_ID~26_combout ;
wire \RegDat2_ID~31_combout ;
wire \always1~1_combout ;
wire \Result_EX~0_combout ;
wire \always1~0_combout ;
wire \Memwrite_EX~0_combout ;
wire \RegDst_ID~0_combout ;
wire \MemToReg_ID~0_combout ;
wire \always1~2_combout ;
wire \care_ID~3_combout ;
wire \MemToReg_ID~q ;
wire \MemToReg_EX~0_combout ;
wire \Result_EX~1_combout ;
wire \Result_EX~2_combout ;
wire \Result_EX~3_combout ;
wire \Result_EX~4_combout ;
wire \Result_EX~5_combout ;
wire \Result_EX~6_combout ;
wire \Result_EX~7_combout ;
wire \Result_EX~8_combout ;
wire \Result_EX~9_combout ;
wire \Result_EX~10_combout ;
wire \Result_EX~11_combout ;
wire \Result_EX[10]~feeder_combout ;
wire \Result_EX~12_combout ;
wire \Result_EX~13_combout ;
wire \Result_EX~14_combout ;
wire \Result_EX~15_combout ;
wire \Result_EX~16_combout ;
wire \Result_EX~17_combout ;
wire \Result_EX~18_combout ;
wire \Result_EX[19]~feeder_combout ;
wire \Result_EX~19_combout ;
wire \Result_EX~20_combout ;
wire \Result_EX~21_combout ;
wire \Result_EX~22_combout ;
wire \Result_EX~23_combout ;
wire \Result_EX~24_combout ;
wire \Result_EX~25_combout ;
wire \Result_EX[24]~feeder_combout ;
wire \Result_EX~26_combout ;
wire \Result_EX~27_combout ;
wire \Result_EX~28_combout ;
wire \Result_EX~29_combout ;
wire \Result_EX~30_combout ;
wire \Result_EX~31_combout ;
wire \halt_ID~0_combout ;
wire \halt_ID~1_combout ;
wire \halt_ID~q ;
wire \halt_EX~0_combout ;
wire \halt_EX~q ;
wire \care_ID~0_combout ;
wire \care_ID~1_combout ;
wire \care_ID~2_combout ;
wire \ALUOP_ID~0_combout ;
wire \ALUOP_ID~1_combout ;
wire \ALUOP_ID~2_combout ;
wire \ALUOP_ID~3_combout ;
wire \ALUOP_ID~4_combout ;
wire \ALUOP_ID~5_combout ;
wire \ALUOP_ID~6_combout ;
wire \ALUOP_ID~7_combout ;
wire \ALUOP_ID~8_combout ;
wire \ALUOP_ID~10_combout ;
wire \ALUOP_ID~9_combout ;
wire \ALUOP_ID~11_combout ;
wire \jump_ID~5_combout ;
wire \RegDst_ID~2_combout ;
wire \RegDst_ID~1_combout ;
wire \RegDst_EX~0_combout ;
wire \RegDst_EX~1_combout ;
wire \RegDst_EX~2_combout ;
wire \RegDst_EX~3_combout ;
wire \RegDst_EX~4_combout ;
wire \RegDst_EX~5_combout ;
wire \RegWen_ID~2_combout ;
wire \RegWen_ID~q ;
wire \RegWen_EX~0_combout ;
wire \RegDst_EX~6_combout ;
wire \RegDst_EX~7_combout ;
wire \RegDst_EX~8_combout ;
wire \RegDst_EX~9_combout ;
wire \Instr_ID~0_combout ;
wire \hazard_Reg_ID~0_combout ;
wire \Instr_ID~1_combout ;
wire \Instr_ID~2_combout ;
wire \Instr_ID~3_combout ;
wire \Memwrite_ID~0_combout ;
wire \Instr_ID~4_combout ;
wire \MemToReg_MEM~feeder_combout ;
wire \Equal3~0_combout ;
wire \ALUSrc2_ID~1_combout ;
wire \ALUSrc2_ID~0_combout ;
wire \ALUSrc2_ID~2_combout ;
wire \ALUSrc2_ID[31]~3_combout ;
wire \Instr_ID~5_combout ;
wire \Instr_ID~6_combout ;
wire \Instr_ID~7_combout ;
wire \Instr_ID~8_combout ;
wire \Instr_ID~9_combout ;
wire \ALUSrc1_ID~0_combout ;
wire \ALUSrc1_ID~1_combout ;
wire \ALUSrc1_ID~2_combout ;
wire \ALUSrc1_ID[31]~3_combout ;
wire \ALUOP_ID~14_combout ;
wire \ALUOP_ID~12_combout ;
wire \ALUOP_ID~13_combout ;
wire \ALUOP_ID~15_combout ;
wire \ALUOP_ID~16_combout ;
wire \ALUSrc1_ID~4_combout ;
wire \ALUSrc1_ID~5_combout ;
wire \ReadData_MEM[30]~feeder_combout ;
wire \Instr_IF~17_combout ;
wire \ALUSrc2_ID~4_combout ;
wire \ALUSrc2_ID~5_combout ;
wire \ALUSrc2_ID~6_combout ;
wire \ALUSrc1_ID~6_combout ;
wire \ALUSrc1_ID~7_combout ;
wire \CalcData_MEM[29]~feeder_combout ;
wire \Instr_IF~24_combout ;
wire \ALUSrc2_ID~7_combout ;
wire \ALUSrc2_ID~8_combout ;
wire \ALUSrc2_ID~9_combout ;
wire \ALUSrc1_ID~8_combout ;
wire \ALUSrc1_ID~9_combout ;
wire \Instr_IF~25_combout ;
wire \ALUSrc2_ID~10_combout ;
wire \ALUSrc2_ID~11_combout ;
wire \ALUSrc2_ID~12_combout ;
wire \ALUSrc1_ID~10_combout ;
wire \ALUSrc1_ID~11_combout ;
wire \ReadData_MEM[27]~feeder_combout ;
wire \Instr_IF~26_combout ;
wire \ALUSrc2_ID~13_combout ;
wire \ALUSrc2_ID~14_combout ;
wire \ALUSrc2_ID~15_combout ;
wire \ALUSrc1_ID~12_combout ;
wire \ALUSrc1_ID~13_combout ;
wire \CalcData_MEM[26]~feeder_combout ;
wire \ALUSrc2_ID~16_combout ;
wire \ALUSrc2_ID~17_combout ;
wire \ALUSrc2_ID~18_combout ;
wire \ALUSrc1_ID~14_combout ;
wire \ALUSrc1_ID~15_combout ;
wire \ReadData_MEM[25]~feeder_combout ;
wire \ALUSrc2_ID~19_combout ;
wire \ALUSrc2_ID~20_combout ;
wire \ALUSrc2_ID~21_combout ;
wire \ALUSrc1_ID~16_combout ;
wire \ALUSrc1_ID~17_combout ;
wire \ALUSrc2_ID~22_combout ;
wire \ALUSrc2_ID~23_combout ;
wire \ALUSrc2_ID~24_combout ;
wire \ALUSrc1_ID~18_combout ;
wire \ALUSrc1_ID~19_combout ;
wire \ALUSrc2_ID~25_combout ;
wire \ALUSrc2_ID~26_combout ;
wire \ALUSrc2_ID~27_combout ;
wire \ALUSrc1_ID~20_combout ;
wire \ALUSrc1_ID~21_combout ;
wire \ReadData_MEM[22]~feeder_combout ;
wire \CalcData_MEM[22]~feeder_combout ;
wire \ALUSrc2_ID~28_combout ;
wire \ALUSrc2_ID~29_combout ;
wire \ALUSrc2_ID~30_combout ;
wire \ALUSrc1_ID~22_combout ;
wire \ALUSrc1_ID~23_combout ;
wire \ReadData_MEM[21]~feeder_combout ;
wire \CalcData_MEM[21]~feeder_combout ;
wire \ALUSrc2_ID~31_combout ;
wire \ALUSrc2_ID~32_combout ;
wire \ALUSrc2_ID~33_combout ;
wire \ALUSrc1_ID~24_combout ;
wire \ALUSrc1_ID~25_combout ;
wire \ReadData_MEM[20]~feeder_combout ;
wire \ALUSrc2_ID~34_combout ;
wire \ALUSrc2_ID~35_combout ;
wire \ALUSrc2_ID~36_combout ;
wire \ALUSrc1_ID~26_combout ;
wire \ALUSrc1_ID~27_combout ;
wire \ALUSrc2_ID~37_combout ;
wire \ALUSrc2_ID~38_combout ;
wire \ALUSrc2_ID~39_combout ;
wire \ALUSrc1_ID~28_combout ;
wire \ALUSrc1_ID~29_combout ;
wire \ReadData_MEM[18]~feeder_combout ;
wire \ALUSrc2_ID~40_combout ;
wire \ALUSrc2_ID~41_combout ;
wire \ALUSrc2_ID~42_combout ;
wire \ALUSrc1_ID~30_combout ;
wire \ALUSrc1_ID~31_combout ;
wire \ALUSrc2_ID~43_combout ;
wire \ALUSrc2_ID~44_combout ;
wire \ALUSrc2_ID~45_combout ;
wire \ALUSrc1_ID~32_combout ;
wire \ALUSrc1_ID~33_combout ;
wire \ReadData_MEM[16]~feeder_combout ;
wire \CalcData_MEM[16]~feeder_combout ;
wire \ALUSrc2_ID~46_combout ;
wire \ALUSrc2_ID~47_combout ;
wire \ALUSrc2_ID~48_combout ;
wire \ALUSrc1_ID~34_combout ;
wire \ALUSrc1_ID~35_combout ;
wire \CalcData_MEM[15]~feeder_combout ;
wire \ALUSrc2_ID~49_combout ;
wire \ALUSrc2_ID~50_combout ;
wire \ALUSrc2_ID~51_combout ;
wire \ALUSrc1_ID~36_combout ;
wire \ALUSrc1_ID~37_combout ;
wire \ReadData_MEM[14]~feeder_combout ;
wire \Instr_IF~23_combout ;
wire \ALUSrc2_ID~52_combout ;
wire \ALUSrc2_ID~53_combout ;
wire \ALUSrc2_ID~54_combout ;
wire \ALUSrc2_ID~55_combout ;
wire \ALUSrc1_ID~38_combout ;
wire \ALUSrc1_ID~39_combout ;
wire \ALUSrc2_ID~56_combout ;
wire \ALUSrc2_ID~57_combout ;
wire \ALUSrc1_ID~40_combout ;
wire \ALUSrc1_ID~41_combout ;
wire \CalcData_MEM[11]~feeder_combout ;
wire \ALUSrc2_ID~58_combout ;
wire \ALUSrc2_ID~59_combout ;
wire \ALUSrc1_ID~42_combout ;
wire \ALUSrc1_ID~43_combout ;
wire \ReadData_MEM[10]~feeder_combout ;
wire \ALUSrc2_ID~60_combout ;
wire \ALUSrc2_ID~61_combout ;
wire \ALUSrc1_ID~44_combout ;
wire \ALUSrc1_ID~45_combout ;
wire \ReadData_MEM[9]~feeder_combout ;
wire \CalcData_MEM[9]~feeder_combout ;
wire \ALUSrc2_ID~62_combout ;
wire \ALUSrc2_ID~63_combout ;
wire \ALUSrc1_ID~46_combout ;
wire \ALUSrc1_ID~47_combout ;
wire \ReadData_MEM[8]~feeder_combout ;
wire \ALUSrc2_ID~64_combout ;
wire \ALUSrc2_ID~65_combout ;
wire \ALUSrc1_ID~48_combout ;
wire \ALUSrc1_ID~49_combout ;
wire \CalcData_MEM[7]~feeder_combout ;
wire \ALUSrc2_ID~66_combout ;
wire \ALUSrc2_ID~67_combout ;
wire \ALUSrc1_ID~50_combout ;
wire \ALUSrc1_ID~51_combout ;
wire \ALUSrc2_ID~68_combout ;
wire \ALUSrc2_ID~69_combout ;
wire \ALUSrc1_ID~52_combout ;
wire \ALUSrc1_ID~53_combout ;
wire \ALUSrc2_ID~70_combout ;
wire \ALUSrc2_ID~71_combout ;
wire \ALUSrc1_ID~54_combout ;
wire \ALUSrc1_ID~55_combout ;
wire \ReadData_MEM[4]~feeder_combout ;
wire \ALUSrc2_ID~72_combout ;
wire \ALUSrc1_ID~56_combout ;
wire \ALUSrc1_ID~57_combout ;
wire \ALUSrc2_ID~73_combout ;
wire \ALUSrc1_ID~58_combout ;
wire \ALUSrc1_ID~59_combout ;
wire \ALUSrc2_ID~74_combout ;
wire \ALUSrc1_ID~60_combout ;
wire \ALUSrc1_ID~61_combout ;
wire \ReadData_MEM[1]~feeder_combout ;
wire \ALUSrc2_ID~75_combout ;
wire \ALUSrc1_ID~62_combout ;
wire \ALUSrc1_ID~63_combout ;
wire \ALUSrc2_ID~76_combout ;
wire \ALUSrc1_ID~64_combout ;
wire \ALUSrc1_ID~65_combout ;
wire \Wdata_EX~1_combout ;
wire \Wdata_EX~0_combout ;
wire \Wdata_EX~2_combout ;
wire \nextPC_IF~0_combout ;
wire \nextPC_ID~0_combout ;
wire \jump_ID~0_combout ;
wire \jump_ID~1_combout ;
wire \jump_ID~2_combout ;
wire \jump_ID~3_combout ;
wire \jump_ID~4_combout ;
wire \nextPC_IF~1_combout ;
wire \nextPC_ID~1_combout ;
wire \nextPC_IF~2_combout ;
wire \nextPC_ID~2_combout ;
wire \Instr_ID~10_combout ;
wire \nextPC_IF~3_combout ;
wire \nextPC_ID~3_combout ;
wire \Instr_ID~11_combout ;
wire \nextPC_IF~4_combout ;
wire \nextPC_ID~4_combout ;
wire \Instr_ID~12_combout ;
wire \nextPC_IF~5_combout ;
wire \nextPC_ID~5_combout ;
wire \Instr_ID~13_combout ;
wire \nextPC_IF~6_combout ;
wire \nextPC_ID~6_combout ;
wire \Instr_ID~14_combout ;
wire \nextPC_IF~7_combout ;
wire \nextPC_ID~7_combout ;
wire \Instr_ID~15_combout ;
wire \nextPC_IF~8_combout ;
wire \nextPC_ID~8_combout ;
wire \Instr_ID~16_combout ;
wire \nextPC_IF~9_combout ;
wire \nextPC_ID~9_combout ;
wire \Instr_ID~17_combout ;
wire \nextPC_IF~10_combout ;
wire \nextPC_ID~10_combout ;
wire \Instr_ID~18_combout ;
wire \nextPC_IF~11_combout ;
wire \nextPC_ID~11_combout ;
wire \Instr_ID~19_combout ;
wire \nextPC_IF~12_combout ;
wire \nextPC_ID~12_combout ;
wire \Instr_ID~20_combout ;
wire \nextPC_IF~13_combout ;
wire \nextPC_ID~13_combout ;
wire \Instr_ID~21_combout ;
wire \nextPC_IF~14_combout ;
wire \nextPC_ID~14_combout ;
wire \Instr_ID~22_combout ;
wire \nextPC_IF~15_combout ;
wire \nextPC_ID~15_combout ;
wire \Instr_ID~23_combout ;
wire \nextPC_IF~16_combout ;
wire \nextPC_ID~16_combout ;
wire \Instr_ID~24_combout ;
wire \nextPC_IF~17_combout ;
wire \nextPC_ID~17_combout ;
wire \Instr_ID~25_combout ;
wire \nextPC_IF~18_combout ;
wire \nextPC_ID~18_combout ;
wire \nextPC_IF~19_combout ;
wire \nextPC_ID~19_combout ;
wire \nextPC_IF~20_combout ;
wire \nextPC_ID~20_combout ;
wire \nextPC_IF~21_combout ;
wire \nextPC_ID~21_combout ;
wire \nextPC_IF~22_combout ;
wire \nextPC_ID~22_combout ;
wire \nextPC_IF~23_combout ;
wire \nextPC_ID~23_combout ;
wire \nextPC_IF~24_combout ;
wire \nextPC_ID~24_combout ;
wire \nextPC_IF~25_combout ;
wire \nextPC_ID~25_combout ;
wire \nextPC_IF~26_combout ;
wire \nextPC_ID~26_combout ;
wire \nextPC_IF~27_combout ;
wire \nextPC_ID~27_combout ;
wire \nextPC_IF~28_combout ;
wire \nextPC_ID~28_combout ;
wire \nextPC_IF~29_combout ;
wire \nextPC_ID~29_combout ;
wire \nextPC_IF~30_combout ;
wire \nextPC_ID~30_combout ;
wire \nextPC_IF~31_combout ;
wire \nextPC_ID~31_combout ;
wire \RegDat2_ID~1_combout ;
wire \Wdata_EX~3_combout ;
wire \Wdata_EX~4_combout ;
wire \RegDat2_ID~2_combout ;
wire \Wdata_EX~5_combout ;
wire \Wdata_EX~6_combout ;
wire \Wdata_EX~7_combout ;
wire \Wdata_EX~8_combout ;
wire \Wdata_EX~9_combout ;
wire \Wdata_EX~10_combout ;
wire \RegDat2_ID~5_combout ;
wire \Wdata_EX~11_combout ;
wire \Wdata_EX~12_combout ;
wire \RegDat2_ID~6_combout ;
wire \Wdata_EX~13_combout ;
wire \Wdata_EX~14_combout ;
wire \RegDat2_ID~7_combout ;
wire \Wdata_EX~15_combout ;
wire \Wdata_EX~16_combout ;
wire \RegDat2_ID~8_combout ;
wire \Wdata_EX~17_combout ;
wire \Wdata_EX~18_combout ;
wire \RegDat2_ID~9_combout ;
wire \Wdata_EX~19_combout ;
wire \Wdata_EX~20_combout ;
wire \RegDat2_ID~10_combout ;
wire \Wdata_EX~21_combout ;
wire \Wdata_EX~22_combout ;
wire \RegDat2_ID~11_combout ;
wire \Wdata_EX~23_combout ;
wire \Wdata_EX~24_combout ;
wire \RegDat2_ID~12_combout ;
wire \Wdata_EX~25_combout ;
wire \Wdata_EX~26_combout ;
wire \Wdata_EX~27_combout ;
wire \Wdata_EX~28_combout ;
wire \RegDat2_ID~14_combout ;
wire \Wdata_EX~29_combout ;
wire \Wdata_EX~30_combout ;
wire \RegDat2_ID~15_combout ;
wire \Wdata_EX~31_combout ;
wire \Wdata_EX~32_combout ;
wire \RegDat2_ID~16_combout ;
wire \Wdata_EX~33_combout ;
wire \Wdata_EX~34_combout ;
wire \Wdata_EX~35_combout ;
wire \Wdata_EX~36_combout ;
wire \RegDat2_ID~18_combout ;
wire \Wdata_EX~37_combout ;
wire \Wdata_EX~38_combout ;
wire \RegDat2_ID~19_combout ;
wire \Wdata_EX~39_combout ;
wire \Wdata_EX~40_combout ;
wire \RegDat2_ID~20_combout ;
wire \Wdata_EX~41_combout ;
wire \Wdata_EX~42_combout ;
wire \RegDat2_ID~21_combout ;
wire \Wdata_EX~43_combout ;
wire \Wdata_EX~44_combout ;
wire \Wdata_EX~45_combout ;
wire \Wdata_EX~46_combout ;
wire \RegDat2_ID~23_combout ;
wire \Wdata_EX~47_combout ;
wire \Wdata_EX~48_combout ;
wire \RegDat2_ID~24_combout ;
wire \Wdata_EX~49_combout ;
wire \Wdata_EX~50_combout ;
wire \RegDat2_ID~25_combout ;
wire \Wdata_EX~51_combout ;
wire \Wdata_EX~52_combout ;
wire \Wdata_EX~53_combout ;
wire \Wdata_EX~54_combout ;
wire \RegDat2_ID~27_combout ;
wire \Wdata_EX~55_combout ;
wire \Wdata_EX~56_combout ;
wire \RegDat2_ID~28_combout ;
wire \Wdata_EX~57_combout ;
wire \Wdata_EX~58_combout ;
wire \RegDat2_ID~29_combout ;
wire \Wdata_EX~59_combout ;
wire \Wdata_EX~60_combout ;
wire \RegDat2_ID~30_combout ;
wire \Wdata_EX~61_combout ;
wire \Wdata_EX~62_combout ;
wire \Wdata_EX~63_combout ;
wire \Wdata_EX~64_combout ;
wire \Instr_IF~0_combout ;
wire \Instr_IF~1_combout ;
wire \Instr_IF~2_combout ;
wire \Instr_IF~3_combout ;
wire \Instr_IF~4_combout ;
wire \Instr_IF~5_combout ;
wire \Instr_IF~6_combout ;
wire \Instr_IF~7_combout ;
wire \Instr_IF~8_combout ;
wire \Instr_IF~9_combout ;
wire \Instr_IF~10_combout ;
wire \Instr_IF~11_combout ;
wire \Instr_IF~12_combout ;
wire \Instr_IF~13_combout ;
wire \Instr_IF~14_combout ;
wire \Instr_IF~15_combout ;
wire \Instr_IF~16_combout ;
wire \Instr_IF~18_combout ;
wire \Instr_IF~19_combout ;
wire \Instr_IF~20_combout ;
wire \Instr_IF~21_combout ;
wire \Instr_IF~22_combout ;
wire \Instr_IF~27_combout ;
wire \Instr_IF~28_combout ;
wire \Instr_IF~29_combout ;
wire \Instr_IF~30_combout ;
wire \Instr_IF~31_combout ;
wire [31:0] nextPC_IF;
wire [1:0] RegDst_ID;
wire [31:0] RegDat2_ID;
wire [31:0] Instr_IF;


// Location: FF_X54_Y32_N11
dffeas \RegDat2_ID[0] (
	.clk(CLK),
	.d(\RegDat2_ID~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[0]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[0] .is_wysiwyg = "true";
defparam \RegDat2_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N21
dffeas \RegDat2_ID[3] (
	.clk(CLK),
	.d(\RegDat2_ID~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[3]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[3] .is_wysiwyg = "true";
defparam \RegDat2_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N19
dffeas \RegDat2_ID[4] (
	.clk(CLK),
	.d(\RegDat2_ID~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[4]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[4] .is_wysiwyg = "true";
defparam \RegDat2_ID[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N7
dffeas \RegDat2_ID[13] (
	.clk(CLK),
	.d(\RegDat2_ID~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[13]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[13] .is_wysiwyg = "true";
defparam \RegDat2_ID[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N17
dffeas \RegDat2_ID[17] (
	.clk(CLK),
	.d(\RegDat2_ID~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[17]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[17] .is_wysiwyg = "true";
defparam \RegDat2_ID[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N3
dffeas \RegDat2_ID[22] (
	.clk(CLK),
	.d(\RegDat2_ID~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[22]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[22] .is_wysiwyg = "true";
defparam \RegDat2_ID[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N23
dffeas \RegDat2_ID[26] (
	.clk(CLK),
	.d(\RegDat2_ID~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[26]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[26] .is_wysiwyg = "true";
defparam \RegDat2_ID[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N7
dffeas \RegDat2_ID[31] (
	.clk(CLK),
	.d(\RegDat2_ID~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[31]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[31] .is_wysiwyg = "true";
defparam \RegDat2_ID[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N4
cycloneive_lcell_comb \RegWen_ID~0 (
// Equation(s):
// \RegWen_ID~0_combout  = (Instr_IF_29 & ((Instr_IF_28) # ((!Instr_IF_31) # (!Instr_IF_26)))) # (!Instr_IF_29 & (!Instr_IF_28 & (Instr_IF_26)))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_28),
	.datac(Instr_IF_26),
	.datad(Instr_IF_31),
	.cin(gnd),
	.combout(\RegWen_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegWen_ID~0 .lut_mask = 16'h9ABA;
defparam \RegWen_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N30
cycloneive_lcell_comb \RegWen_ID~1 (
// Equation(s):
// \RegWen_ID~1_combout  = (Instr_IF_30 & (!Decoder0 & ((!Selector11)))) # (!Instr_IF_30 & ((\RegWen_ID~0_combout ) # ((!Decoder0 & !Selector11))))

	.dataa(Instr_IF_30),
	.datab(Decoder0),
	.datac(\RegWen_ID~0_combout ),
	.datad(Selector111),
	.cin(gnd),
	.combout(\RegWen_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegWen_ID~1 .lut_mask = 16'h5073;
defparam \RegWen_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \RegDat2_ID~0 (
// Equation(s):
// \RegDat2_ID~0_combout  = (rfifrdat2_0 & !\branch~0_combout )

	.dataa(rfifrdat2_0),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~0 .lut_mask = 16'h00AA;
defparam \RegDat2_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \RegDat2_ID~3 (
// Equation(s):
// \RegDat2_ID~3_combout  = (!\branch~0_combout  & rfifrdat2_3)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_3),
	.cin(gnd),
	.combout(\RegDat2_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~3 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \RegDat2_ID~4 (
// Equation(s):
// \RegDat2_ID~4_combout  = (rfifrdat2_4 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_4),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDat2_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~4 .lut_mask = 16'h0C0C;
defparam \RegDat2_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \RegDat2_ID~13 (
// Equation(s):
// \RegDat2_ID~13_combout  = (rfifrdat2_13 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_13),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~13 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \RegDat2_ID~17 (
// Equation(s):
// \RegDat2_ID~17_combout  = (rfifrdat2_17 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_17),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~17_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~17 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \RegDat2_ID~22 (
// Equation(s):
// \RegDat2_ID~22_combout  = (rfifrdat2_22 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(rfifrdat2_22),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~22_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~22 .lut_mask = 16'h00F0;
defparam \RegDat2_ID~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \RegDat2_ID~26 (
// Equation(s):
// \RegDat2_ID~26_combout  = (rfifrdat2_26 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_26),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~26_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~26 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \RegDat2_ID~31 (
// Equation(s):
// \RegDat2_ID~31_combout  = (rfifrdat2_31 & !\branch~0_combout )

	.dataa(rfifrdat2_31),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~31_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~31 .lut_mask = 16'h00AA;
defparam \RegDat2_ID~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N17
dffeas \Result_EX[1] (
	.clk(CLK),
	.d(\Result_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_1),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[1] .is_wysiwyg = "true";
defparam \Result_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas Memwrite_EX(
	.clk(CLK),
	.d(gnd),
	.asdata(\Memwrite_EX~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Memwrite_EX1),
	.prn(vcc));
// synopsys translate_off
defparam Memwrite_EX.is_wysiwyg = "true";
defparam Memwrite_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N17
dffeas MemToReg_EX(
	.clk(CLK),
	.d(gnd),
	.asdata(\MemToReg_EX~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(MemToReg_EX1),
	.prn(vcc));
// synopsys translate_off
defparam MemToReg_EX.is_wysiwyg = "true";
defparam MemToReg_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N15
dffeas \Result_EX[0] (
	.clk(CLK),
	.d(\Result_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_0),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[0] .is_wysiwyg = "true";
defparam \Result_EX[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N21
dffeas \Result_EX[3] (
	.clk(CLK),
	.d(\Result_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_3),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[3] .is_wysiwyg = "true";
defparam \Result_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N27
dffeas \Result_EX[2] (
	.clk(CLK),
	.d(\Result_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_2),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[2] .is_wysiwyg = "true";
defparam \Result_EX[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N1
dffeas \Result_EX[5] (
	.clk(CLK),
	.d(\Result_EX~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_5),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[5] .is_wysiwyg = "true";
defparam \Result_EX[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N25
dffeas \Result_EX[4] (
	.clk(CLK),
	.d(\Result_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_4),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[4] .is_wysiwyg = "true";
defparam \Result_EX[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N13
dffeas \Result_EX[7] (
	.clk(CLK),
	.d(\Result_EX~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_7),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[7] .is_wysiwyg = "true";
defparam \Result_EX[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N7
dffeas \Result_EX[6] (
	.clk(CLK),
	.d(\Result_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_6),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[6] .is_wysiwyg = "true";
defparam \Result_EX[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N5
dffeas \Result_EX[9] (
	.clk(CLK),
	.d(\Result_EX~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_9),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[9] .is_wysiwyg = "true";
defparam \Result_EX[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N27
dffeas \Result_EX[8] (
	.clk(CLK),
	.d(\Result_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_8),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[8] .is_wysiwyg = "true";
defparam \Result_EX[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N21
dffeas \Result_EX[11] (
	.clk(CLK),
	.d(\Result_EX~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_11),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[11] .is_wysiwyg = "true";
defparam \Result_EX[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N1
dffeas \Result_EX[10] (
	.clk(CLK),
	.d(\Result_EX[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_10),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[10] .is_wysiwyg = "true";
defparam \Result_EX[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N5
dffeas \Result_EX[13] (
	.clk(CLK),
	.d(\Result_EX~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_13),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[13] .is_wysiwyg = "true";
defparam \Result_EX[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N29
dffeas \Result_EX[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Result_EX~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_12),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[12] .is_wysiwyg = "true";
defparam \Result_EX[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N19
dffeas \Result_EX[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Result_EX~14_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_15),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[15] .is_wysiwyg = "true";
defparam \Result_EX[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N31
dffeas \Result_EX[14] (
	.clk(CLK),
	.d(\Result_EX~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_14),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[14] .is_wysiwyg = "true";
defparam \Result_EX[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N17
dffeas \Result_EX[17] (
	.clk(CLK),
	.d(\Result_EX~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_17),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[17] .is_wysiwyg = "true";
defparam \Result_EX[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N7
dffeas \Result_EX[16] (
	.clk(CLK),
	.d(\Result_EX~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_16),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[16] .is_wysiwyg = "true";
defparam \Result_EX[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N21
dffeas \Result_EX[19] (
	.clk(CLK),
	.d(\Result_EX[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_19),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[19] .is_wysiwyg = "true";
defparam \Result_EX[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N15
dffeas \Result_EX[18] (
	.clk(CLK),
	.d(\Result_EX~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_18),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[18] .is_wysiwyg = "true";
defparam \Result_EX[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N7
dffeas \Result_EX[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Result_EX~20_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_21),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[21] .is_wysiwyg = "true";
defparam \Result_EX[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \Result_EX[20] (
	.clk(CLK),
	.d(\Result_EX~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_20),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[20] .is_wysiwyg = "true";
defparam \Result_EX[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N25
dffeas \Result_EX[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Result_EX~22_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_23),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[23] .is_wysiwyg = "true";
defparam \Result_EX[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N17
dffeas \Result_EX[22] (
	.clk(CLK),
	.d(\Result_EX~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_22),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[22] .is_wysiwyg = "true";
defparam \Result_EX[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \Result_EX[25] (
	.clk(CLK),
	.d(\Result_EX~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_25),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[25] .is_wysiwyg = "true";
defparam \Result_EX[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N13
dffeas \Result_EX[24] (
	.clk(CLK),
	.d(\Result_EX[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_24),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[24] .is_wysiwyg = "true";
defparam \Result_EX[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N31
dffeas \Result_EX[27] (
	.clk(CLK),
	.d(\Result_EX~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_27),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[27] .is_wysiwyg = "true";
defparam \Result_EX[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N21
dffeas \Result_EX[26] (
	.clk(CLK),
	.d(\Result_EX~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_26),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[26] .is_wysiwyg = "true";
defparam \Result_EX[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \Result_EX[29] (
	.clk(CLK),
	.d(\Result_EX~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_29),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[29] .is_wysiwyg = "true";
defparam \Result_EX[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N1
dffeas \Result_EX[28] (
	.clk(CLK),
	.d(\Result_EX~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_28),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[28] .is_wysiwyg = "true";
defparam \Result_EX[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N15
dffeas \Result_EX[31] (
	.clk(CLK),
	.d(\Result_EX~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_31),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[31] .is_wysiwyg = "true";
defparam \Result_EX[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N11
dffeas \Result_EX[30] (
	.clk(CLK),
	.d(\Result_EX~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Result_EX_30),
	.prn(vcc));
// synopsys translate_off
defparam \Result_EX[30] .is_wysiwyg = "true";
defparam \Result_EX[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N23
dffeas halt_MEM(
	.clk(CLK),
	.d(gnd),
	.asdata(\halt_EX~q ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(halt_MEM1),
	.prn(vcc));
// synopsys translate_off
defparam halt_MEM.is_wysiwyg = "true";
defparam halt_MEM.power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N29
dffeas care_ID(
	.clk(CLK),
	.d(\care_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(care_ID1),
	.prn(vcc));
// synopsys translate_off
defparam care_ID.is_wysiwyg = "true";
defparam care_ID.power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N25
dffeas \ALUOP_ID[1] (
	.clk(CLK),
	.d(\ALUOP_ID~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOP_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOP_ID[1] .is_wysiwyg = "true";
defparam \ALUOP_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N3
dffeas \ALUOP_ID[3] (
	.clk(CLK),
	.d(\ALUOP_ID~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOP_ID_3),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOP_ID[3] .is_wysiwyg = "true";
defparam \ALUOP_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N27
dffeas \ALUOP_ID[2] (
	.clk(CLK),
	.d(\ALUOP_ID~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOP_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOP_ID[2] .is_wysiwyg = "true";
defparam \ALUOP_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \RegDst_EX[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\RegDst_EX~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_EX_0),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_EX[0] .is_wysiwyg = "true";
defparam \RegDst_EX[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N21
dffeas \RegDst_EX[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\RegDst_EX~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_EX_1),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_EX[1] .is_wysiwyg = "true";
defparam \RegDst_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N7
dffeas \RegDst_EX[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\RegDst_EX~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_EX_2),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_EX[2] .is_wysiwyg = "true";
defparam \RegDst_EX[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N15
dffeas RegWen_EX(
	.clk(CLK),
	.d(gnd),
	.asdata(\RegWen_EX~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegWen_EX1),
	.prn(vcc));
// synopsys translate_off
defparam RegWen_EX.is_wysiwyg = "true";
defparam RegWen_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N5
dffeas \RegDst_EX[3] (
	.clk(CLK),
	.d(\RegDst_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_EX_3),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_EX[3] .is_wysiwyg = "true";
defparam \RegDst_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N27
dffeas \RegDst_EX[4] (
	.clk(CLK),
	.d(\RegDst_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_EX_4),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_EX[4] .is_wysiwyg = "true";
defparam \RegDst_EX[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N23
dffeas \Instr_ID[16] (
	.clk(CLK),
	.d(\Instr_ID~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_16),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[16] .is_wysiwyg = "true";
defparam \Instr_ID[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N23
dffeas hazard_Reg_ID(
	.clk(CLK),
	.d(gnd),
	.asdata(\hazard_Reg_ID~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(hazard_Reg_ID1),
	.prn(vcc));
// synopsys translate_off
defparam hazard_Reg_ID.is_wysiwyg = "true";
defparam hazard_Reg_ID.power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N7
dffeas \Instr_ID[17] (
	.clk(CLK),
	.d(\Instr_ID~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_17),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[17] .is_wysiwyg = "true";
defparam \Instr_ID[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N31
dffeas \Instr_ID[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Instr_ID~2_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_18),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[18] .is_wysiwyg = "true";
defparam \Instr_ID[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N27
dffeas \Instr_ID[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Instr_ID~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_19),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[19] .is_wysiwyg = "true";
defparam \Instr_ID[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N25
dffeas Memwrite_ID(
	.clk(CLK),
	.d(gnd),
	.asdata(\Memwrite_ID~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Memwrite_ID1),
	.prn(vcc));
// synopsys translate_off
defparam Memwrite_ID.is_wysiwyg = "true";
defparam Memwrite_ID.power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \Instr_ID[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Instr_ID~4_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_20),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[20] .is_wysiwyg = "true";
defparam \Instr_ID[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N17
dffeas \ReadData_MEM[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_31),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[31] .is_wysiwyg = "true";
defparam \ReadData_MEM[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N7
dffeas \CalcData_MEM[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_31),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[31] .is_wysiwyg = "true";
defparam \CalcData_MEM[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas MemToReg_MEM(
	.clk(CLK),
	.d(\MemToReg_MEM~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(MemToReg_MEM1),
	.prn(vcc));
// synopsys translate_off
defparam MemToReg_MEM.is_wysiwyg = "true";
defparam MemToReg_MEM.power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N17
dffeas RegWen_MEM(
	.clk(CLK),
	.d(gnd),
	.asdata(RegWen_EX1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegWen_MEM1),
	.prn(vcc));
// synopsys translate_off
defparam RegWen_MEM.is_wysiwyg = "true";
defparam RegWen_MEM.power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \RegDst_MEM[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(RegDst_EX_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_MEM_0),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_MEM[0] .is_wysiwyg = "true";
defparam \RegDst_MEM[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N23
dffeas \RegDst_MEM[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(RegDst_EX_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_MEM_1),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_MEM[1] .is_wysiwyg = "true";
defparam \RegDst_MEM[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N31
dffeas \RegDst_MEM[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(RegDst_EX_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_MEM_4),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_MEM[4] .is_wysiwyg = "true";
defparam \RegDst_MEM[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \RegDst_MEM[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(RegDst_EX_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_MEM_3),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_MEM[3] .is_wysiwyg = "true";
defparam \RegDst_MEM[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \RegDst_MEM[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(RegDst_EX_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_MEM_2),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_MEM[2] .is_wysiwyg = "true";
defparam \RegDst_MEM[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \ALUSrc2_ID[31] (
	.clk(CLK),
	.d(\ALUSrc2_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_31),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[31] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N21
dffeas \Instr_ID[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Instr_ID~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_21),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[21] .is_wysiwyg = "true";
defparam \Instr_ID[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N21
dffeas \Instr_ID[22] (
	.clk(CLK),
	.d(\Instr_ID~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_22),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[22] .is_wysiwyg = "true";
defparam \Instr_ID[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N17
dffeas \Instr_ID[24] (
	.clk(CLK),
	.d(\Instr_ID~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_24),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[24] .is_wysiwyg = "true";
defparam \Instr_ID[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N17
dffeas \Instr_ID[25] (
	.clk(CLK),
	.d(\Instr_ID~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_25),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[25] .is_wysiwyg = "true";
defparam \Instr_ID[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N25
dffeas \Instr_ID[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Instr_ID~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_23),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[23] .is_wysiwyg = "true";
defparam \Instr_ID[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N13
dffeas \ALUSrc1_ID[31] (
	.clk(CLK),
	.d(\ALUSrc1_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_31),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[31] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N7
dffeas \ALUOP_ID[0] (
	.clk(CLK),
	.d(\ALUOP_ID~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOP_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOP_ID[0] .is_wysiwyg = "true";
defparam \ALUOP_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N29
dffeas \ALUSrc1_ID[30] (
	.clk(CLK),
	.d(\ALUSrc1_ID~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_30),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[30] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N19
dffeas \ReadData_MEM[30] (
	.clk(CLK),
	.d(\ReadData_MEM[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_30),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[30] .is_wysiwyg = "true";
defparam \ReadData_MEM[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N13
dffeas \CalcData_MEM[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_30),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[30] .is_wysiwyg = "true";
defparam \CalcData_MEM[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N29
dffeas \ALUSrc2_ID[30] (
	.clk(CLK),
	.d(\ALUSrc2_ID~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_30),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[30] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N9
dffeas \ALUSrc1_ID[29] (
	.clk(CLK),
	.d(\ALUSrc1_ID~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_29),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[29] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N7
dffeas \ReadData_MEM[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_29),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[29] .is_wysiwyg = "true";
defparam \ReadData_MEM[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N3
dffeas \CalcData_MEM[29] (
	.clk(CLK),
	.d(\CalcData_MEM[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_29),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[29] .is_wysiwyg = "true";
defparam \CalcData_MEM[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N13
dffeas \ALUSrc2_ID[29] (
	.clk(CLK),
	.d(\ALUSrc2_ID~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_29),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[29] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N7
dffeas \ALUSrc1_ID[28] (
	.clk(CLK),
	.d(\ALUSrc1_ID~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_28),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[28] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N27
dffeas \ReadData_MEM[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_28),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[28] .is_wysiwyg = "true";
defparam \ReadData_MEM[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N5
dffeas \CalcData_MEM[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_28),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[28] .is_wysiwyg = "true";
defparam \CalcData_MEM[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N3
dffeas \ALUSrc2_ID[28] (
	.clk(CLK),
	.d(\ALUSrc2_ID~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_28),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[28] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N25
dffeas \ALUSrc1_ID[27] (
	.clk(CLK),
	.d(\ALUSrc1_ID~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_27),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[27] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N19
dffeas \ReadData_MEM[27] (
	.clk(CLK),
	.d(\ReadData_MEM[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_27),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[27] .is_wysiwyg = "true";
defparam \ReadData_MEM[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N29
dffeas \CalcData_MEM[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_27),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[27] .is_wysiwyg = "true";
defparam \CalcData_MEM[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N15
dffeas \ALUSrc2_ID[27] (
	.clk(CLK),
	.d(\ALUSrc2_ID~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_27),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[27] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N15
dffeas \ALUSrc1_ID[26] (
	.clk(CLK),
	.d(\ALUSrc1_ID~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_26),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[26] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N3
dffeas \ReadData_MEM[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_26),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[26] .is_wysiwyg = "true";
defparam \ReadData_MEM[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N5
dffeas \CalcData_MEM[26] (
	.clk(CLK),
	.d(\CalcData_MEM[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_26),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[26] .is_wysiwyg = "true";
defparam \CalcData_MEM[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N15
dffeas \ALUSrc2_ID[26] (
	.clk(CLK),
	.d(\ALUSrc2_ID~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_26),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[26] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N29
dffeas \ALUSrc1_ID[25] (
	.clk(CLK),
	.d(\ALUSrc1_ID~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_25),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[25] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N27
dffeas \ReadData_MEM[25] (
	.clk(CLK),
	.d(\ReadData_MEM[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_25),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[25] .is_wysiwyg = "true";
defparam \ReadData_MEM[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N29
dffeas \CalcData_MEM[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_25),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[25] .is_wysiwyg = "true";
defparam \CalcData_MEM[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N17
dffeas \ALUSrc2_ID[25] (
	.clk(CLK),
	.d(\ALUSrc2_ID~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_25),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[25] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N29
dffeas \ALUSrc1_ID[24] (
	.clk(CLK),
	.d(\ALUSrc1_ID~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_24),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[24] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \ReadData_MEM[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_24),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[24] .is_wysiwyg = "true";
defparam \ReadData_MEM[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N17
dffeas \CalcData_MEM[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_24),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[24] .is_wysiwyg = "true";
defparam \CalcData_MEM[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N21
dffeas \ALUSrc2_ID[24] (
	.clk(CLK),
	.d(\ALUSrc2_ID~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_24),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[24] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N31
dffeas \ALUSrc1_ID[23] (
	.clk(CLK),
	.d(\ALUSrc1_ID~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_23),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[23] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N7
dffeas \ReadData_MEM[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_23),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[23] .is_wysiwyg = "true";
defparam \ReadData_MEM[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N25
dffeas \CalcData_MEM[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_23),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[23] .is_wysiwyg = "true";
defparam \CalcData_MEM[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N23
dffeas \ALUSrc2_ID[23] (
	.clk(CLK),
	.d(\ALUSrc2_ID~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_23),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[23] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N1
dffeas \ALUSrc1_ID[22] (
	.clk(CLK),
	.d(\ALUSrc1_ID~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_22),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[22] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N17
dffeas \ReadData_MEM[22] (
	.clk(CLK),
	.d(\ReadData_MEM[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_22),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[22] .is_wysiwyg = "true";
defparam \ReadData_MEM[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N15
dffeas \CalcData_MEM[22] (
	.clk(CLK),
	.d(\CalcData_MEM[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_22),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[22] .is_wysiwyg = "true";
defparam \CalcData_MEM[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N27
dffeas \ALUSrc2_ID[22] (
	.clk(CLK),
	.d(\ALUSrc2_ID~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_22),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[22] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N23
dffeas \ALUSrc1_ID[21] (
	.clk(CLK),
	.d(\ALUSrc1_ID~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_21),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[21] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N5
dffeas \ReadData_MEM[21] (
	.clk(CLK),
	.d(\ReadData_MEM[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_21),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[21] .is_wysiwyg = "true";
defparam \ReadData_MEM[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N11
dffeas \CalcData_MEM[21] (
	.clk(CLK),
	.d(\CalcData_MEM[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_21),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[21] .is_wysiwyg = "true";
defparam \CalcData_MEM[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N29
dffeas \ALUSrc2_ID[21] (
	.clk(CLK),
	.d(\ALUSrc2_ID~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_21),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[21] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \ALUSrc1_ID[20] (
	.clk(CLK),
	.d(\ALUSrc1_ID~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_20),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[20] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N29
dffeas \ReadData_MEM[20] (
	.clk(CLK),
	.d(\ReadData_MEM[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_20),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[20] .is_wysiwyg = "true";
defparam \ReadData_MEM[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N11
dffeas \CalcData_MEM[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_20),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[20] .is_wysiwyg = "true";
defparam \CalcData_MEM[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N27
dffeas \ALUSrc2_ID[20] (
	.clk(CLK),
	.d(\ALUSrc2_ID~36_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_20),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[20] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N5
dffeas \ALUSrc1_ID[19] (
	.clk(CLK),
	.d(\ALUSrc1_ID~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_19),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[19] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N29
dffeas \ReadData_MEM[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_19),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[19] .is_wysiwyg = "true";
defparam \ReadData_MEM[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \CalcData_MEM[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_19),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[19] .is_wysiwyg = "true";
defparam \CalcData_MEM[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N17
dffeas \ALUSrc2_ID[19] (
	.clk(CLK),
	.d(\ALUSrc2_ID~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_19),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[19] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N23
dffeas \ALUSrc1_ID[18] (
	.clk(CLK),
	.d(\ALUSrc1_ID~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_18),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[18] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N9
dffeas \ReadData_MEM[18] (
	.clk(CLK),
	.d(\ReadData_MEM[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_18),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[18] .is_wysiwyg = "true";
defparam \ReadData_MEM[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N27
dffeas \CalcData_MEM[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_18),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[18] .is_wysiwyg = "true";
defparam \CalcData_MEM[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N13
dffeas \ALUSrc2_ID[18] (
	.clk(CLK),
	.d(\ALUSrc2_ID~42_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_18),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[18] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \ALUSrc1_ID[17] (
	.clk(CLK),
	.d(\ALUSrc1_ID~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_17),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[17] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N5
dffeas \ReadData_MEM[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_17),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[17] .is_wysiwyg = "true";
defparam \ReadData_MEM[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N13
dffeas \CalcData_MEM[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_17),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[17] .is_wysiwyg = "true";
defparam \CalcData_MEM[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N31
dffeas \ALUSrc2_ID[17] (
	.clk(CLK),
	.d(\ALUSrc2_ID~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_17),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[17] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N21
dffeas \ALUSrc1_ID[16] (
	.clk(CLK),
	.d(\ALUSrc1_ID~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_16),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[16] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N29
dffeas \ReadData_MEM[16] (
	.clk(CLK),
	.d(\ReadData_MEM[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_16),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[16] .is_wysiwyg = "true";
defparam \ReadData_MEM[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N21
dffeas \CalcData_MEM[16] (
	.clk(CLK),
	.d(\CalcData_MEM[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_16),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[16] .is_wysiwyg = "true";
defparam \CalcData_MEM[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N3
dffeas \ALUSrc2_ID[16] (
	.clk(CLK),
	.d(\ALUSrc2_ID~48_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_16),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[16] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \ALUSrc1_ID[15] (
	.clk(CLK),
	.d(\ALUSrc1_ID~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_15),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[15] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N3
dffeas \ReadData_MEM[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_15),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[15] .is_wysiwyg = "true";
defparam \ReadData_MEM[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N21
dffeas \CalcData_MEM[15] (
	.clk(CLK),
	.d(\CalcData_MEM[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_15),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[15] .is_wysiwyg = "true";
defparam \CalcData_MEM[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N31
dffeas \ALUSrc2_ID[15] (
	.clk(CLK),
	.d(\ALUSrc2_ID~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_15),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[15] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \ALUSrc1_ID[14] (
	.clk(CLK),
	.d(\ALUSrc1_ID~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_14),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[14] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N27
dffeas \ReadData_MEM[14] (
	.clk(CLK),
	.d(\ReadData_MEM[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_14),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[14] .is_wysiwyg = "true";
defparam \ReadData_MEM[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N9
dffeas \CalcData_MEM[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_14),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[14] .is_wysiwyg = "true";
defparam \CalcData_MEM[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N1
dffeas \ALUSrc2_ID[14] (
	.clk(CLK),
	.d(\ALUSrc2_ID~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_14),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[14] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N1
dffeas \ReadData_MEM[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_13),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[13] .is_wysiwyg = "true";
defparam \ReadData_MEM[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N31
dffeas \CalcData_MEM[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_13),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[13] .is_wysiwyg = "true";
defparam \CalcData_MEM[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N29
dffeas \ALUSrc2_ID[13] (
	.clk(CLK),
	.d(\ALUSrc2_ID~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_13),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[13] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N17
dffeas \ALUSrc1_ID[13] (
	.clk(CLK),
	.d(\ALUSrc1_ID~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_13),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[13] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N29
dffeas \ReadData_MEM[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_12),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[12] .is_wysiwyg = "true";
defparam \ReadData_MEM[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N23
dffeas \CalcData_MEM[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_12),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[12] .is_wysiwyg = "true";
defparam \CalcData_MEM[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N5
dffeas \ALUSrc2_ID[12] (
	.clk(CLK),
	.d(\ALUSrc2_ID~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_12),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[12] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N15
dffeas \ALUSrc1_ID[12] (
	.clk(CLK),
	.d(\ALUSrc1_ID~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_12),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[12] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y30_N23
dffeas \ReadData_MEM[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_11),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[11] .is_wysiwyg = "true";
defparam \ReadData_MEM[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y30_N25
dffeas \CalcData_MEM[11] (
	.clk(CLK),
	.d(\CalcData_MEM[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_11),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[11] .is_wysiwyg = "true";
defparam \CalcData_MEM[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N31
dffeas \ALUSrc2_ID[11] (
	.clk(CLK),
	.d(\ALUSrc2_ID~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_11),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[11] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N21
dffeas \ALUSrc1_ID[11] (
	.clk(CLK),
	.d(\ALUSrc1_ID~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_11),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[11] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y30_N29
dffeas \ReadData_MEM[10] (
	.clk(CLK),
	.d(\ReadData_MEM[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_10),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[10] .is_wysiwyg = "true";
defparam \ReadData_MEM[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y30_N3
dffeas \CalcData_MEM[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_10),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[10] .is_wysiwyg = "true";
defparam \CalcData_MEM[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N17
dffeas \ALUSrc2_ID[10] (
	.clk(CLK),
	.d(\ALUSrc2_ID~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_10),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[10] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N29
dffeas \ALUSrc1_ID[10] (
	.clk(CLK),
	.d(\ALUSrc1_ID~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_10),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[10] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N27
dffeas \ReadData_MEM[9] (
	.clk(CLK),
	.d(\ReadData_MEM[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_9),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[9] .is_wysiwyg = "true";
defparam \ReadData_MEM[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N9
dffeas \CalcData_MEM[9] (
	.clk(CLK),
	.d(\CalcData_MEM[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_9),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[9] .is_wysiwyg = "true";
defparam \CalcData_MEM[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N21
dffeas \ALUSrc2_ID[9] (
	.clk(CLK),
	.d(\ALUSrc2_ID~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_9),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[9] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N11
dffeas \ALUSrc1_ID[9] (
	.clk(CLK),
	.d(\ALUSrc1_ID~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_9),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[9] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \ReadData_MEM[8] (
	.clk(CLK),
	.d(\ReadData_MEM[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_8),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[8] .is_wysiwyg = "true";
defparam \ReadData_MEM[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N19
dffeas \CalcData_MEM[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_8),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[8] .is_wysiwyg = "true";
defparam \CalcData_MEM[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N13
dffeas \ALUSrc2_ID[8] (
	.clk(CLK),
	.d(\ALUSrc2_ID~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_8),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[8] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \ALUSrc1_ID[8] (
	.clk(CLK),
	.d(\ALUSrc1_ID~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_8),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[8] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N11
dffeas \ReadData_MEM[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_7),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[7] .is_wysiwyg = "true";
defparam \ReadData_MEM[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N1
dffeas \CalcData_MEM[7] (
	.clk(CLK),
	.d(\CalcData_MEM[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_7),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[7] .is_wysiwyg = "true";
defparam \CalcData_MEM[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \ALUSrc2_ID[7] (
	.clk(CLK),
	.d(\ALUSrc2_ID~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_7),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[7] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N9
dffeas \ALUSrc1_ID[7] (
	.clk(CLK),
	.d(\ALUSrc1_ID~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_7),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[7] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N23
dffeas \ReadData_MEM[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_6),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[6] .is_wysiwyg = "true";
defparam \ReadData_MEM[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N13
dffeas \CalcData_MEM[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_6),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[6] .is_wysiwyg = "true";
defparam \CalcData_MEM[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N9
dffeas \ALUSrc2_ID[6] (
	.clk(CLK),
	.d(\ALUSrc2_ID~69_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_6),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[6] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N21
dffeas \ALUSrc1_ID[6] (
	.clk(CLK),
	.d(\ALUSrc1_ID~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_6),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[6] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N15
dffeas \ReadData_MEM[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_5),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[5] .is_wysiwyg = "true";
defparam \ReadData_MEM[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N5
dffeas \CalcData_MEM[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_5),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[5] .is_wysiwyg = "true";
defparam \CalcData_MEM[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \ALUSrc2_ID[5] (
	.clk(CLK),
	.d(\ALUSrc2_ID~71_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_5),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[5] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N11
dffeas \ALUSrc1_ID[5] (
	.clk(CLK),
	.d(\ALUSrc1_ID~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_5),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[5] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N29
dffeas \ReadData_MEM[4] (
	.clk(CLK),
	.d(\ReadData_MEM[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_4),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[4] .is_wysiwyg = "true";
defparam \ReadData_MEM[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N23
dffeas \CalcData_MEM[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_4),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[4] .is_wysiwyg = "true";
defparam \CalcData_MEM[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N3
dffeas \ALUSrc2_ID[4] (
	.clk(CLK),
	.d(\ALUSrc2_ID~72_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_4),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[4] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N13
dffeas \ALUSrc1_ID[4] (
	.clk(CLK),
	.d(\ALUSrc1_ID~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_4),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[4] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N5
dffeas \ReadData_MEM[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_3),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[3] .is_wysiwyg = "true";
defparam \ReadData_MEM[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N3
dffeas \CalcData_MEM[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_3),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[3] .is_wysiwyg = "true";
defparam \CalcData_MEM[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \ALUSrc2_ID[3] (
	.clk(CLK),
	.d(\ALUSrc2_ID~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_3),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[3] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N1
dffeas \ALUSrc1_ID[3] (
	.clk(CLK),
	.d(\ALUSrc1_ID~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_3),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[3] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N3
dffeas \ReadData_MEM[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_2),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[2] .is_wysiwyg = "true";
defparam \ReadData_MEM[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N23
dffeas \CalcData_MEM[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_2),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[2] .is_wysiwyg = "true";
defparam \CalcData_MEM[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N11
dffeas \ALUSrc2_ID[2] (
	.clk(CLK),
	.d(\ALUSrc2_ID~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[2] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N19
dffeas \ALUSrc1_ID[2] (
	.clk(CLK),
	.d(\ALUSrc1_ID~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[2] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N25
dffeas \ReadData_MEM[1] (
	.clk(CLK),
	.d(\ReadData_MEM[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_1),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[1] .is_wysiwyg = "true";
defparam \ReadData_MEM[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N7
dffeas \CalcData_MEM[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_1),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[1] .is_wysiwyg = "true";
defparam \CalcData_MEM[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N15
dffeas \ALUSrc2_ID[1] (
	.clk(CLK),
	.d(\ALUSrc2_ID~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[1] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N7
dffeas \ALUSrc1_ID[1] (
	.clk(CLK),
	.d(\ALUSrc1_ID~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[1] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N25
dffeas \ReadData_MEM[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ReadData_MEM_0),
	.prn(vcc));
// synopsys translate_off
defparam \ReadData_MEM[0] .is_wysiwyg = "true";
defparam \ReadData_MEM[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N11
dffeas \CalcData_MEM[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(Result_EX_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(CalcData_MEM_0),
	.prn(vcc));
// synopsys translate_off
defparam \CalcData_MEM[0] .is_wysiwyg = "true";
defparam \CalcData_MEM[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \ALUSrc2_ID[0] (
	.clk(CLK),
	.d(\ALUSrc2_ID~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc2_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc2_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc2_ID[0] .is_wysiwyg = "true";
defparam \ALUSrc2_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N27
dffeas \ALUSrc1_ID[0] (
	.clk(CLK),
	.d(\ALUSrc1_ID~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc1_ID[31]~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUSrc1_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \ALUSrc1_ID[0] .is_wysiwyg = "true";
defparam \ALUSrc1_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N5
dffeas \Wdata_EX[0] (
	.clk(CLK),
	.d(\Wdata_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_0),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[0] .is_wysiwyg = "true";
defparam \Wdata_EX[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N7
dffeas \nextPC_ID[1] (
	.clk(CLK),
	.d(\nextPC_ID~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[1] .is_wysiwyg = "true";
defparam \nextPC_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N9
dffeas \jump_ID[0] (
	.clk(CLK),
	.d(\jump_ID~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(jump_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \jump_ID[0] .is_wysiwyg = "true";
defparam \jump_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N29
dffeas \jump_ID[1] (
	.clk(CLK),
	.d(\jump_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(jump_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \jump_ID[1] .is_wysiwyg = "true";
defparam \jump_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N11
dffeas \jump_ID[2] (
	.clk(CLK),
	.d(\jump_ID~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(jump_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \jump_ID[2] .is_wysiwyg = "true";
defparam \jump_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N13
dffeas \nextPC_ID[0] (
	.clk(CLK),
	.d(\nextPC_ID~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[0] .is_wysiwyg = "true";
defparam \nextPC_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N19
dffeas \nextPC_ID[3] (
	.clk(CLK),
	.d(\nextPC_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_3),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[3] .is_wysiwyg = "true";
defparam \nextPC_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N1
dffeas \Instr_ID[1] (
	.clk(CLK),
	.d(\Instr_ID~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_1),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[1] .is_wysiwyg = "true";
defparam \Instr_ID[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N29
dffeas \nextPC_ID[2] (
	.clk(CLK),
	.d(\nextPC_ID~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[2] .is_wysiwyg = "true";
defparam \nextPC_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N3
dffeas \Instr_ID[0] (
	.clk(CLK),
	.d(\Instr_ID~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_0),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[0] .is_wysiwyg = "true";
defparam \Instr_ID[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N9
dffeas \nextPC_ID[5] (
	.clk(CLK),
	.d(\nextPC_ID~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_5),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[5] .is_wysiwyg = "true";
defparam \nextPC_ID[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N11
dffeas \Instr_ID[3] (
	.clk(CLK),
	.d(\Instr_ID~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_3),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[3] .is_wysiwyg = "true";
defparam \Instr_ID[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N5
dffeas \nextPC_ID[4] (
	.clk(CLK),
	.d(\nextPC_ID~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_4),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[4] .is_wysiwyg = "true";
defparam \nextPC_ID[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N25
dffeas \Instr_ID[2] (
	.clk(CLK),
	.d(\Instr_ID~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_2),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[2] .is_wysiwyg = "true";
defparam \Instr_ID[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N13
dffeas \nextPC_ID[7] (
	.clk(CLK),
	.d(\nextPC_ID~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_7),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[7] .is_wysiwyg = "true";
defparam \nextPC_ID[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N17
dffeas \Instr_ID[5] (
	.clk(CLK),
	.d(\Instr_ID~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_5),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[5] .is_wysiwyg = "true";
defparam \Instr_ID[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N11
dffeas \nextPC_ID[6] (
	.clk(CLK),
	.d(\nextPC_ID~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_6),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[6] .is_wysiwyg = "true";
defparam \nextPC_ID[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N23
dffeas \Instr_ID[4] (
	.clk(CLK),
	.d(\Instr_ID~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_4),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[4] .is_wysiwyg = "true";
defparam \Instr_ID[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N15
dffeas \nextPC_ID[9] (
	.clk(CLK),
	.d(\nextPC_ID~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_9),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[9] .is_wysiwyg = "true";
defparam \nextPC_ID[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N21
dffeas \Instr_ID[7] (
	.clk(CLK),
	.d(\Instr_ID~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_7),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[7] .is_wysiwyg = "true";
defparam \Instr_ID[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N11
dffeas \nextPC_ID[8] (
	.clk(CLK),
	.d(\nextPC_ID~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_8),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[8] .is_wysiwyg = "true";
defparam \nextPC_ID[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N25
dffeas \Instr_ID[6] (
	.clk(CLK),
	.d(\Instr_ID~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_6),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[6] .is_wysiwyg = "true";
defparam \Instr_ID[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N29
dffeas \nextPC_ID[11] (
	.clk(CLK),
	.d(\nextPC_ID~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_11),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[11] .is_wysiwyg = "true";
defparam \nextPC_ID[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N31
dffeas \Instr_ID[9] (
	.clk(CLK),
	.d(\Instr_ID~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_9),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[9] .is_wysiwyg = "true";
defparam \Instr_ID[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N15
dffeas \nextPC_ID[10] (
	.clk(CLK),
	.d(\nextPC_ID~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_10),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[10] .is_wysiwyg = "true";
defparam \nextPC_ID[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N1
dffeas \Instr_ID[8] (
	.clk(CLK),
	.d(\Instr_ID~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_8),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[8] .is_wysiwyg = "true";
defparam \Instr_ID[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N7
dffeas \nextPC_ID[13] (
	.clk(CLK),
	.d(\nextPC_ID~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_13),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[13] .is_wysiwyg = "true";
defparam \nextPC_ID[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N15
dffeas \Instr_ID[11] (
	.clk(CLK),
	.d(\Instr_ID~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_11),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[11] .is_wysiwyg = "true";
defparam \Instr_ID[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N31
dffeas \nextPC_ID[12] (
	.clk(CLK),
	.d(\nextPC_ID~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_12),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[12] .is_wysiwyg = "true";
defparam \nextPC_ID[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N11
dffeas \Instr_ID[10] (
	.clk(CLK),
	.d(\Instr_ID~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_10),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[10] .is_wysiwyg = "true";
defparam \Instr_ID[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N9
dffeas \nextPC_ID[15] (
	.clk(CLK),
	.d(\nextPC_ID~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_15),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[15] .is_wysiwyg = "true";
defparam \nextPC_ID[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N13
dffeas \Instr_ID[13] (
	.clk(CLK),
	.d(\Instr_ID~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_13),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[13] .is_wysiwyg = "true";
defparam \Instr_ID[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N27
dffeas \nextPC_ID[14] (
	.clk(CLK),
	.d(\nextPC_ID~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_14),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[14] .is_wysiwyg = "true";
defparam \nextPC_ID[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N31
dffeas \Instr_ID[12] (
	.clk(CLK),
	.d(\Instr_ID~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_12),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[12] .is_wysiwyg = "true";
defparam \Instr_ID[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N5
dffeas \nextPC_ID[17] (
	.clk(CLK),
	.d(\nextPC_ID~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_17),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[17] .is_wysiwyg = "true";
defparam \nextPC_ID[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N15
dffeas \Instr_ID[15] (
	.clk(CLK),
	.d(\Instr_ID~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_15),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[15] .is_wysiwyg = "true";
defparam \Instr_ID[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N31
dffeas \nextPC_ID[16] (
	.clk(CLK),
	.d(\nextPC_ID~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_16),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[16] .is_wysiwyg = "true";
defparam \nextPC_ID[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N25
dffeas \Instr_ID[14] (
	.clk(CLK),
	.d(\Instr_ID~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_ID_14),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_ID[14] .is_wysiwyg = "true";
defparam \Instr_ID[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N7
dffeas \nextPC_ID[19] (
	.clk(CLK),
	.d(\nextPC_ID~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_19),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[19] .is_wysiwyg = "true";
defparam \nextPC_ID[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N25
dffeas \nextPC_ID[18] (
	.clk(CLK),
	.d(\nextPC_ID~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_18),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[18] .is_wysiwyg = "true";
defparam \nextPC_ID[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N7
dffeas \nextPC_ID[21] (
	.clk(CLK),
	.d(\nextPC_ID~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_21),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[21] .is_wysiwyg = "true";
defparam \nextPC_ID[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N29
dffeas \nextPC_ID[20] (
	.clk(CLK),
	.d(\nextPC_ID~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_20),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[20] .is_wysiwyg = "true";
defparam \nextPC_ID[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N31
dffeas \nextPC_ID[23] (
	.clk(CLK),
	.d(\nextPC_ID~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_23),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[23] .is_wysiwyg = "true";
defparam \nextPC_ID[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N17
dffeas \nextPC_ID[22] (
	.clk(CLK),
	.d(\nextPC_ID~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_22),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[22] .is_wysiwyg = "true";
defparam \nextPC_ID[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N5
dffeas \nextPC_ID[25] (
	.clk(CLK),
	.d(\nextPC_ID~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_25),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[25] .is_wysiwyg = "true";
defparam \nextPC_ID[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N17
dffeas \nextPC_ID[24] (
	.clk(CLK),
	.d(\nextPC_ID~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_24),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[24] .is_wysiwyg = "true";
defparam \nextPC_ID[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N9
dffeas \nextPC_ID[27] (
	.clk(CLK),
	.d(\nextPC_ID~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_27),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[27] .is_wysiwyg = "true";
defparam \nextPC_ID[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N11
dffeas \nextPC_ID[26] (
	.clk(CLK),
	.d(\nextPC_ID~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_26),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[26] .is_wysiwyg = "true";
defparam \nextPC_ID[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N21
dffeas \nextPC_ID[29] (
	.clk(CLK),
	.d(\nextPC_ID~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_29),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[29] .is_wysiwyg = "true";
defparam \nextPC_ID[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N31
dffeas \nextPC_ID[28] (
	.clk(CLK),
	.d(\nextPC_ID~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_28),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[28] .is_wysiwyg = "true";
defparam \nextPC_ID[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N25
dffeas \nextPC_ID[31] (
	.clk(CLK),
	.d(\nextPC_ID~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_31),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[31] .is_wysiwyg = "true";
defparam \nextPC_ID[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N19
dffeas \nextPC_ID[30] (
	.clk(CLK),
	.d(\nextPC_ID~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_ID_30),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_ID[30] .is_wysiwyg = "true";
defparam \nextPC_ID[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas \Wdata_EX[1] (
	.clk(CLK),
	.d(\Wdata_EX~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_1),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[1] .is_wysiwyg = "true";
defparam \Wdata_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N25
dffeas \Wdata_EX[2] (
	.clk(CLK),
	.d(\Wdata_EX~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_2),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[2] .is_wysiwyg = "true";
defparam \Wdata_EX[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N15
dffeas \Wdata_EX[3] (
	.clk(CLK),
	.d(\Wdata_EX~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_3),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[3] .is_wysiwyg = "true";
defparam \Wdata_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N9
dffeas \Wdata_EX[4] (
	.clk(CLK),
	.d(\Wdata_EX~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_4),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[4] .is_wysiwyg = "true";
defparam \Wdata_EX[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N21
dffeas \Wdata_EX[5] (
	.clk(CLK),
	.d(\Wdata_EX~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_5),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[5] .is_wysiwyg = "true";
defparam \Wdata_EX[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N11
dffeas \Wdata_EX[6] (
	.clk(CLK),
	.d(\Wdata_EX~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_6),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[6] .is_wysiwyg = "true";
defparam \Wdata_EX[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N5
dffeas \Wdata_EX[7] (
	.clk(CLK),
	.d(\Wdata_EX~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_7),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[7] .is_wysiwyg = "true";
defparam \Wdata_EX[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N29
dffeas \Wdata_EX[8] (
	.clk(CLK),
	.d(\Wdata_EX~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_8),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[8] .is_wysiwyg = "true";
defparam \Wdata_EX[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N13
dffeas \Wdata_EX[9] (
	.clk(CLK),
	.d(\Wdata_EX~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_9),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[9] .is_wysiwyg = "true";
defparam \Wdata_EX[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N1
dffeas \Wdata_EX[10] (
	.clk(CLK),
	.d(\Wdata_EX~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_10),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[10] .is_wysiwyg = "true";
defparam \Wdata_EX[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N5
dffeas \Wdata_EX[11] (
	.clk(CLK),
	.d(\Wdata_EX~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_11),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[11] .is_wysiwyg = "true";
defparam \Wdata_EX[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \Wdata_EX[12] (
	.clk(CLK),
	.d(\Wdata_EX~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_12),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[12] .is_wysiwyg = "true";
defparam \Wdata_EX[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N17
dffeas \Wdata_EX[13] (
	.clk(CLK),
	.d(\Wdata_EX~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_13),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[13] .is_wysiwyg = "true";
defparam \Wdata_EX[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N25
dffeas \Wdata_EX[14] (
	.clk(CLK),
	.d(\Wdata_EX~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_14),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[14] .is_wysiwyg = "true";
defparam \Wdata_EX[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N3
dffeas \Wdata_EX[15] (
	.clk(CLK),
	.d(\Wdata_EX~32_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_15),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[15] .is_wysiwyg = "true";
defparam \Wdata_EX[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N21
dffeas \Wdata_EX[16] (
	.clk(CLK),
	.d(\Wdata_EX~34_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_16),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[16] .is_wysiwyg = "true";
defparam \Wdata_EX[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N7
dffeas \Wdata_EX[17] (
	.clk(CLK),
	.d(\Wdata_EX~36_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_17),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[17] .is_wysiwyg = "true";
defparam \Wdata_EX[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N9
dffeas \Wdata_EX[18] (
	.clk(CLK),
	.d(\Wdata_EX~38_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_18),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[18] .is_wysiwyg = "true";
defparam \Wdata_EX[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N29
dffeas \Wdata_EX[19] (
	.clk(CLK),
	.d(\Wdata_EX~40_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_19),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[19] .is_wysiwyg = "true";
defparam \Wdata_EX[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N7
dffeas \Wdata_EX[20] (
	.clk(CLK),
	.d(\Wdata_EX~42_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_20),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[20] .is_wysiwyg = "true";
defparam \Wdata_EX[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N27
dffeas \Wdata_EX[21] (
	.clk(CLK),
	.d(\Wdata_EX~44_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_21),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[21] .is_wysiwyg = "true";
defparam \Wdata_EX[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \Wdata_EX[22] (
	.clk(CLK),
	.d(\Wdata_EX~46_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_22),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[22] .is_wysiwyg = "true";
defparam \Wdata_EX[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N29
dffeas \Wdata_EX[23] (
	.clk(CLK),
	.d(\Wdata_EX~48_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_23),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[23] .is_wysiwyg = "true";
defparam \Wdata_EX[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \Wdata_EX[24] (
	.clk(CLK),
	.d(\Wdata_EX~50_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_24),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[24] .is_wysiwyg = "true";
defparam \Wdata_EX[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N11
dffeas \Wdata_EX[25] (
	.clk(CLK),
	.d(\Wdata_EX~52_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_25),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[25] .is_wysiwyg = "true";
defparam \Wdata_EX[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N19
dffeas \Wdata_EX[26] (
	.clk(CLK),
	.d(\Wdata_EX~54_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_26),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[26] .is_wysiwyg = "true";
defparam \Wdata_EX[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N15
dffeas \Wdata_EX[27] (
	.clk(CLK),
	.d(\Wdata_EX~56_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_27),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[27] .is_wysiwyg = "true";
defparam \Wdata_EX[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N31
dffeas \Wdata_EX[28] (
	.clk(CLK),
	.d(\Wdata_EX~58_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_28),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[28] .is_wysiwyg = "true";
defparam \Wdata_EX[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N9
dffeas \Wdata_EX[29] (
	.clk(CLK),
	.d(\Wdata_EX~60_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_29),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[29] .is_wysiwyg = "true";
defparam \Wdata_EX[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N7
dffeas \Wdata_EX[30] (
	.clk(CLK),
	.d(\Wdata_EX~62_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_30),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[30] .is_wysiwyg = "true";
defparam \Wdata_EX[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N21
dffeas \Wdata_EX[31] (
	.clk(CLK),
	.d(\Wdata_EX~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Wdata_EX_31),
	.prn(vcc));
// synopsys translate_off
defparam \Wdata_EX[31] .is_wysiwyg = "true";
defparam \Wdata_EX[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N21
dffeas \Instr_IF[30] (
	.clk(CLK),
	.d(\Instr_IF~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_30),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[30] .is_wysiwyg = "true";
defparam \Instr_IF[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N31
dffeas \Instr_IF[28] (
	.clk(CLK),
	.d(\Instr_IF~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_28),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[28] .is_wysiwyg = "true";
defparam \Instr_IF[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N1
dffeas \Instr_IF[26] (
	.clk(CLK),
	.d(\Instr_IF~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_26),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[26] .is_wysiwyg = "true";
defparam \Instr_IF[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N23
dffeas \Instr_IF[27] (
	.clk(CLK),
	.d(\Instr_IF~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_27),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[27] .is_wysiwyg = "true";
defparam \Instr_IF[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N21
dffeas \Instr_IF[29] (
	.clk(CLK),
	.d(\Instr_IF~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_29),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[29] .is_wysiwyg = "true";
defparam \Instr_IF[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N25
dffeas \Instr_IF[5] (
	.clk(CLK),
	.d(\Instr_IF~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_5),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[5] .is_wysiwyg = "true";
defparam \Instr_IF[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N27
dffeas \Instr_IF[4] (
	.clk(CLK),
	.d(\Instr_IF~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_4),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[4] .is_wysiwyg = "true";
defparam \Instr_IF[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N19
dffeas \Instr_IF[2] (
	.clk(CLK),
	.d(\Instr_IF~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_2),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[2] .is_wysiwyg = "true";
defparam \Instr_IF[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N15
dffeas \Instr_IF[3] (
	.clk(CLK),
	.d(\Instr_IF~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_3),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[3] .is_wysiwyg = "true";
defparam \Instr_IF[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N27
dffeas \Instr_IF[0] (
	.clk(CLK),
	.d(\Instr_IF~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_0),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[0] .is_wysiwyg = "true";
defparam \Instr_IF[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \Instr_IF[1] (
	.clk(CLK),
	.d(\Instr_IF~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_1),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[1] .is_wysiwyg = "true";
defparam \Instr_IF[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N15
dffeas \Instr_IF[31] (
	.clk(CLK),
	.d(\Instr_IF~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_31),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[31] .is_wysiwyg = "true";
defparam \Instr_IF[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N1
dffeas \Instr_IF[16] (
	.clk(CLK),
	.d(\Instr_IF~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_16),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[16] .is_wysiwyg = "true";
defparam \Instr_IF[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N21
dffeas \Instr_IF[17] (
	.clk(CLK),
	.d(\Instr_IF~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_17),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[17] .is_wysiwyg = "true";
defparam \Instr_IF[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N19
dffeas \Instr_IF[18] (
	.clk(CLK),
	.d(\Instr_IF~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_18),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[18] .is_wysiwyg = "true";
defparam \Instr_IF[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N31
dffeas \Instr_IF[19] (
	.clk(CLK),
	.d(\Instr_IF~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_19),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[19] .is_wysiwyg = "true";
defparam \Instr_IF[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N5
dffeas \Instr_IF[20] (
	.clk(CLK),
	.d(\Instr_IF~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_20),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[20] .is_wysiwyg = "true";
defparam \Instr_IF[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N1
dffeas \Instr_IF[21] (
	.clk(CLK),
	.d(\Instr_IF~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_21),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[21] .is_wysiwyg = "true";
defparam \Instr_IF[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N27
dffeas \Instr_IF[22] (
	.clk(CLK),
	.d(\Instr_IF~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_22),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[22] .is_wysiwyg = "true";
defparam \Instr_IF[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N5
dffeas \Instr_IF[24] (
	.clk(CLK),
	.d(\Instr_IF~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_24),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[24] .is_wysiwyg = "true";
defparam \Instr_IF[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N7
dffeas \Instr_IF[25] (
	.clk(CLK),
	.d(\Instr_IF~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_25),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[25] .is_wysiwyg = "true";
defparam \Instr_IF[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N13
dffeas \Instr_IF[23] (
	.clk(CLK),
	.d(\Instr_IF~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_23),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[23] .is_wysiwyg = "true";
defparam \Instr_IF[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N31
dffeas \Instr_IF[10] (
	.clk(CLK),
	.d(\Instr_IF~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_10),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[10] .is_wysiwyg = "true";
defparam \Instr_IF[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N27
dffeas \Instr_IF[9] (
	.clk(CLK),
	.d(\Instr_IF~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_9),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[9] .is_wysiwyg = "true";
defparam \Instr_IF[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N5
dffeas \Instr_IF[8] (
	.clk(CLK),
	.d(\Instr_IF~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_8),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[8] .is_wysiwyg = "true";
defparam \Instr_IF[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N25
dffeas \Instr_IF[7] (
	.clk(CLK),
	.d(\Instr_IF~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_7),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[7] .is_wysiwyg = "true";
defparam \Instr_IF[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N7
dffeas \Instr_IF[6] (
	.clk(CLK),
	.d(\Instr_IF~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF_6),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[6] .is_wysiwyg = "true";
defparam \Instr_IF[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// \always1~1_combout  = (\always1~0_combout  & ((!src2_hazard_t1) # (!always01)))

	.dataa(\always1~0_combout ),
	.datab(always0),
	.datac(gnd),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\always1~1_combout ),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'h22AA;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \Result_EX~0 (
// Equation(s):
// \Result_EX~0_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_1)) # (!\Equal8~0_combout  & ((Selector30)))))

	.dataa(\always1~1_combout ),
	.datab(Equal8),
	.datac(nextPC_ID_1),
	.datad(Selector30),
	.cin(gnd),
	.combout(\Result_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~0 .lut_mask = 16'hA280;
defparam \Result_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// \always1~0_combout  = ((!always03 & ((!MemToReg_MEM1) # (!src1_hazard_t)))) # (!MemToReg_EX1)

	.dataa(src1_hazard_t),
	.datab(MemToReg_MEM1),
	.datac(always01),
	.datad(MemToReg_EX1),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h07FF;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \Memwrite_EX~0 (
// Equation(s):
// \Memwrite_EX~0_combout  = (Memwrite_ID1 & (\always1~0_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(Memwrite_ID1),
	.datab(\always1~0_combout ),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Memwrite_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \Memwrite_EX~0 .lut_mask = 16'h0888;
defparam \Memwrite_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N10
cycloneive_lcell_comb \RegDst_ID~0 (
// Equation(s):
// \RegDst_ID~0_combout  = (!Instr_IF_30 & (WideOr21 & !\branch~0_combout ))

	.dataa(Instr_IF_30),
	.datab(gnd),
	.datac(WideOr21),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDst_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_ID~0 .lut_mask = 16'h0050;
defparam \RegDst_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N26
cycloneive_lcell_comb \MemToReg_ID~0 (
// Equation(s):
// \MemToReg_ID~0_combout  = (!Instr_IF_29 & (Instr_IF_31 & \RegDst_ID~0_combout ))

	.dataa(gnd),
	.datab(Instr_IF_29),
	.datac(Instr_IF_31),
	.datad(\RegDst_ID~0_combout ),
	.cin(gnd),
	.combout(\MemToReg_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \MemToReg_ID~0 .lut_mask = 16'h3000;
defparam \MemToReg_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \always1~2 (
// Equation(s):
// \always1~2_combout  = ((always01 & (src2_hazard_t1)) # (!always01 & (!src2_hazard_t1 & src2_hazard_t2))) # (!\always1~0_combout )

	.dataa(always0),
	.datab(\always1~0_combout ),
	.datac(src2_hazard_t),
	.datad(src2_hazard_t1),
	.cin(gnd),
	.combout(\always1~2_combout ),
	.cout());
// synopsys translate_off
defparam \always1~2 .lut_mask = 16'hB7B3;
defparam \always1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \care_ID~3 (
// Equation(s):
// \care_ID~3_combout  = (!\always1~2_combout  & always1)

	.dataa(gnd),
	.datab(\always1~2_combout ),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(\care_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \care_ID~3 .lut_mask = 16'h3030;
defparam \care_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N27
dffeas MemToReg_ID(
	.clk(CLK),
	.d(\MemToReg_ID~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\MemToReg_ID~q ),
	.prn(vcc));
// synopsys translate_off
defparam MemToReg_ID.is_wysiwyg = "true";
defparam MemToReg_ID.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N16
cycloneive_lcell_comb \MemToReg_EX~0 (
// Equation(s):
// \MemToReg_EX~0_combout  = (\MemToReg_ID~q  & (\always1~0_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(\MemToReg_ID~q ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\MemToReg_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \MemToReg_EX~0 .lut_mask = 16'h7000;
defparam \MemToReg_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \Result_EX~1 (
// Equation(s):
// \Result_EX~1_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_0)) # (!\Equal8~0_combout  & ((Selector31)))))

	.dataa(\always1~1_combout ),
	.datab(Equal8),
	.datac(nextPC_ID_0),
	.datad(Selector31),
	.cin(gnd),
	.combout(\Result_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~1 .lut_mask = 16'hA280;
defparam \Result_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \Result_EX~2 (
// Equation(s):
// \Result_EX~2_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_3))) # (!\Equal8~0_combout  & (Selector28))))

	.dataa(\always1~1_combout ),
	.datab(Equal8),
	.datac(Selector28),
	.datad(nextPC_ID_3),
	.cin(gnd),
	.combout(\Result_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~2 .lut_mask = 16'hA820;
defparam \Result_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \Result_EX~3 (
// Equation(s):
// \Result_EX~3_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_2)) # (!\Equal8~0_combout  & ((Selector29)))))

	.dataa(\always1~1_combout ),
	.datab(Equal8),
	.datac(nextPC_ID_2),
	.datad(Selector29),
	.cin(gnd),
	.combout(\Result_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~3 .lut_mask = 16'hA280;
defparam \Result_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \Result_EX~4 (
// Equation(s):
// \Result_EX~4_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_5)) # (!\Equal8~0_combout  & ((Selector26)))))

	.dataa(\always1~1_combout ),
	.datab(Equal8),
	.datac(nextPC_ID_5),
	.datad(Selector26),
	.cin(gnd),
	.combout(\Result_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~4 .lut_mask = 16'hA280;
defparam \Result_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N24
cycloneive_lcell_comb \Result_EX~5 (
// Equation(s):
// \Result_EX~5_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_4)) # (!\Equal8~0_combout  & ((Selector27)))))

	.dataa(nextPC_ID_4),
	.datab(Equal8),
	.datac(\always1~1_combout ),
	.datad(Selector27),
	.cin(gnd),
	.combout(\Result_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~5 .lut_mask = 16'hB080;
defparam \Result_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Result_EX~6 (
// Equation(s):
// \Result_EX~6_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_7)) # (!\Equal8~0_combout  & ((Selector24)))))

	.dataa(nextPC_ID_7),
	.datab(\always1~1_combout ),
	.datac(Selector24),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~6 .lut_mask = 16'h88C0;
defparam \Result_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N6
cycloneive_lcell_comb \Result_EX~7 (
// Equation(s):
// \Result_EX~7_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_6))) # (!\Equal8~0_combout  & (Selector25))))

	.dataa(Selector25),
	.datab(nextPC_ID_6),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~7 .lut_mask = 16'hC0A0;
defparam \Result_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \Result_EX~8 (
// Equation(s):
// \Result_EX~8_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_9)) # (!\Equal8~0_combout  & ((Selector22)))))

	.dataa(nextPC_ID_9),
	.datab(Selector22),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~8 .lut_mask = 16'hA0C0;
defparam \Result_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \Result_EX~9 (
// Equation(s):
// \Result_EX~9_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_8)) # (!\Equal8~0_combout  & ((Selector23)))))

	.dataa(nextPC_ID_8),
	.datab(Selector23),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~9 .lut_mask = 16'hA0C0;
defparam \Result_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \Result_EX~10 (
// Equation(s):
// \Result_EX~10_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_11))) # (!\Equal8~0_combout  & (Selector20))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(Selector20),
	.datad(nextPC_ID_11),
	.cin(gnd),
	.combout(\Result_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~10 .lut_mask = 16'hC840;
defparam \Result_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N20
cycloneive_lcell_comb \Result_EX~11 (
// Equation(s):
// \Result_EX~11_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_10)) # (!\Equal8~0_combout  & ((Selector21)))))

	.dataa(Equal8),
	.datab(nextPC_ID_10),
	.datac(Selector21),
	.datad(\always1~1_combout ),
	.cin(gnd),
	.combout(\Result_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~11 .lut_mask = 16'hD800;
defparam \Result_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \Result_EX[10]~feeder (
// Equation(s):
// \Result_EX[10]~feeder_combout  = \Result_EX~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Result_EX~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Result_EX[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX[10]~feeder .lut_mask = 16'hF0F0;
defparam \Result_EX[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N4
cycloneive_lcell_comb \Result_EX~12 (
// Equation(s):
// \Result_EX~12_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_13)) # (!\Equal8~0_combout  & ((Selector18)))))

	.dataa(\always1~1_combout ),
	.datab(nextPC_ID_13),
	.datac(Selector18),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~12 .lut_mask = 16'h88A0;
defparam \Result_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \Result_EX~13 (
// Equation(s):
// \Result_EX~13_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_12))) # (!\Equal8~0_combout  & (Selector19))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(Selector19),
	.datad(nextPC_ID_12),
	.cin(gnd),
	.combout(\Result_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~13 .lut_mask = 16'hC840;
defparam \Result_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N24
cycloneive_lcell_comb \Result_EX~14 (
// Equation(s):
// \Result_EX~14_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_15)) # (!\Equal8~0_combout  & ((Selector16)))))

	.dataa(\always1~1_combout ),
	.datab(nextPC_ID_15),
	.datac(Equal8),
	.datad(Selector16),
	.cin(gnd),
	.combout(\Result_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~14 .lut_mask = 16'h8A80;
defparam \Result_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N30
cycloneive_lcell_comb \Result_EX~15 (
// Equation(s):
// \Result_EX~15_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_14))) # (!\Equal8~0_combout  & (Selector17))))

	.dataa(Selector17),
	.datab(Equal8),
	.datac(\always1~1_combout ),
	.datad(nextPC_ID_14),
	.cin(gnd),
	.combout(\Result_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~15 .lut_mask = 16'hE020;
defparam \Result_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Result_EX~16 (
// Equation(s):
// \Result_EX~16_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_17)) # (!\Equal8~0_combout  & ((Selector14)))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(nextPC_ID_17),
	.datad(Selector14),
	.cin(gnd),
	.combout(\Result_EX~16_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~16 .lut_mask = 16'hC480;
defparam \Result_EX~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \Result_EX~17 (
// Equation(s):
// \Result_EX~17_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_16))) # (!\Equal8~0_combout  & (Selector15))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(Selector15),
	.datad(nextPC_ID_16),
	.cin(gnd),
	.combout(\Result_EX~17_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~17 .lut_mask = 16'hC840;
defparam \Result_EX~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \Result_EX~18 (
// Equation(s):
// \Result_EX~18_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_19))) # (!\Equal8~0_combout  & (Selector12))))

	.dataa(\always1~1_combout ),
	.datab(Selector12),
	.datac(nextPC_ID_19),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~18_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~18 .lut_mask = 16'hA088;
defparam \Result_EX~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \Result_EX[19]~feeder (
// Equation(s):
// \Result_EX[19]~feeder_combout  = \Result_EX~18_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Result_EX~18_combout ),
	.cin(gnd),
	.combout(\Result_EX[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX[19]~feeder .lut_mask = 16'hFF00;
defparam \Result_EX[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \Result_EX~19 (
// Equation(s):
// \Result_EX~19_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_18)) # (!\Equal8~0_combout  & ((Selector13)))))

	.dataa(Equal8),
	.datab(nextPC_ID_18),
	.datac(Selector13),
	.datad(\always1~1_combout ),
	.cin(gnd),
	.combout(\Result_EX~19_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~19 .lut_mask = 16'hD800;
defparam \Result_EX~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \Result_EX~20 (
// Equation(s):
// \Result_EX~20_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_21)) # (!\Equal8~0_combout  & ((Selector10)))))

	.dataa(Equal8),
	.datab(nextPC_ID_21),
	.datac(Selector10),
	.datad(\always1~1_combout ),
	.cin(gnd),
	.combout(\Result_EX~20_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~20 .lut_mask = 16'hD800;
defparam \Result_EX~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \Result_EX~21 (
// Equation(s):
// \Result_EX~21_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_20))) # (!\Equal8~0_combout  & (Selector11))))

	.dataa(Selector11),
	.datab(nextPC_ID_20),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~21_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~21 .lut_mask = 16'hC0A0;
defparam \Result_EX~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N6
cycloneive_lcell_comb \Result_EX~22 (
// Equation(s):
// \Result_EX~22_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_23)) # (!\Equal8~0_combout  & ((Selector8)))))

	.dataa(\always1~1_combout ),
	.datab(nextPC_ID_23),
	.datac(Equal8),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Result_EX~22_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~22 .lut_mask = 16'h8A80;
defparam \Result_EX~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \Result_EX~23 (
// Equation(s):
// \Result_EX~23_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_22)) # (!\Equal8~0_combout  & ((Selector9)))))

	.dataa(\always1~1_combout ),
	.datab(nextPC_ID_22),
	.datac(Selector9),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~23_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~23 .lut_mask = 16'h88A0;
defparam \Result_EX~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \Result_EX~24 (
// Equation(s):
// \Result_EX~24_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_25))) # (!\Equal8~0_combout  & (Selector6))))

	.dataa(Selector6),
	.datab(nextPC_ID_25),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~24_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~24 .lut_mask = 16'hC0A0;
defparam \Result_EX~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N2
cycloneive_lcell_comb \Result_EX~25 (
// Equation(s):
// \Result_EX~25_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_24))) # (!\Equal8~0_combout  & (Selector7))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(Selector7),
	.datad(nextPC_ID_24),
	.cin(gnd),
	.combout(\Result_EX~25_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~25 .lut_mask = 16'hC840;
defparam \Result_EX~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \Result_EX[24]~feeder (
// Equation(s):
// \Result_EX[24]~feeder_combout  = \Result_EX~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Result_EX~25_combout ),
	.cin(gnd),
	.combout(\Result_EX[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX[24]~feeder .lut_mask = 16'hFF00;
defparam \Result_EX[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \Result_EX~26 (
// Equation(s):
// \Result_EX~26_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_27)) # (!\Equal8~0_combout  & ((Selector4)))))

	.dataa(nextPC_ID_27),
	.datab(Selector4),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~26_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~26 .lut_mask = 16'hA0C0;
defparam \Result_EX~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Result_EX~27 (
// Equation(s):
// \Result_EX~27_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & (nextPC_ID_26)) # (!\Equal8~0_combout  & ((Selector5)))))

	.dataa(nextPC_ID_26),
	.datab(Selector5),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~27_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~27 .lut_mask = 16'hA0C0;
defparam \Result_EX~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Result_EX~28 (
// Equation(s):
// \Result_EX~28_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_29))) # (!\Equal8~0_combout  & (Selector2))))

	.dataa(Selector2),
	.datab(\always1~1_combout ),
	.datac(nextPC_ID_29),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~28_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~28 .lut_mask = 16'hC088;
defparam \Result_EX~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Result_EX~29 (
// Equation(s):
// \Result_EX~29_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_28))) # (!\Equal8~0_combout  & (Selector3))))

	.dataa(Selector3),
	.datab(nextPC_ID_28),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~29_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~29 .lut_mask = 16'hC0A0;
defparam \Result_EX~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \Result_EX~30 (
// Equation(s):
// \Result_EX~30_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_31))) # (!\Equal8~0_combout  & (Selector0))))

	.dataa(Equal8),
	.datab(\always1~1_combout ),
	.datac(Selector0),
	.datad(nextPC_ID_31),
	.cin(gnd),
	.combout(\Result_EX~30_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~30 .lut_mask = 16'hC840;
defparam \Result_EX~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \Result_EX~31 (
// Equation(s):
// \Result_EX~31_combout  = (\always1~1_combout  & ((\Equal8~0_combout  & ((nextPC_ID_30))) # (!\Equal8~0_combout  & (Selector1))))

	.dataa(Selector1),
	.datab(nextPC_ID_30),
	.datac(\always1~1_combout ),
	.datad(Equal8),
	.cin(gnd),
	.combout(\Result_EX~31_combout ),
	.cout());
// synopsys translate_off
defparam \Result_EX~31 .lut_mask = 16'hC0A0;
defparam \Result_EX~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N2
cycloneive_lcell_comb \halt_ID~0 (
// Equation(s):
// \halt_ID~0_combout  = (Instr_IF_30) # ((Instr_IF_31 & ((!WideOr21))) # (!Instr_IF_31 & (WideOr11)))

	.dataa(Instr_IF_30),
	.datab(WideOr11),
	.datac(Instr_IF_31),
	.datad(WideOr21),
	.cin(gnd),
	.combout(\halt_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_ID~0 .lut_mask = 16'hAEFE;
defparam \halt_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N18
cycloneive_lcell_comb \halt_ID~1 (
// Equation(s):
// \halt_ID~1_combout  = (\halt_ID~0_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\halt_ID~0_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\halt_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \halt_ID~1 .lut_mask = 16'h00F0;
defparam \halt_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N19
dffeas halt_ID(
	.clk(CLK),
	.d(\halt_ID~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\halt_ID~q ),
	.prn(vcc));
// synopsys translate_off
defparam halt_ID.is_wysiwyg = "true";
defparam halt_ID.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N8
cycloneive_lcell_comb \halt_EX~0 (
// Equation(s):
// \halt_EX~0_combout  = (\halt_ID~q  & (\always1~0_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(\halt_ID~q ),
	.datac(\always1~0_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(\halt_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_EX~0 .lut_mask = 16'h40C0;
defparam \halt_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N9
dffeas halt_EX(
	.clk(CLK),
	.d(\halt_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\halt_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam halt_EX.is_wysiwyg = "true";
defparam halt_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N0
cycloneive_lcell_comb \care_ID~0 (
// Equation(s):
// \care_ID~0_combout  = (!Instr_IF_3 & (Instr_IF_5 & (!Instr_IF_4 & !Instr_IF_2)))

	.dataa(Instr_IF_3),
	.datab(Instr_IF_5),
	.datac(Instr_IF_4),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(\care_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \care_ID~0 .lut_mask = 16'h0004;
defparam \care_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N18
cycloneive_lcell_comb \care_ID~1 (
// Equation(s):
// \care_ID~1_combout  = (Selector14 & ((Instr_IF_29) # ((\care_ID~0_combout  & !Instr_IF_0))))

	.dataa(Selector141),
	.datab(Instr_IF_29),
	.datac(\care_ID~0_combout ),
	.datad(Instr_IF_0),
	.cin(gnd),
	.combout(\care_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \care_ID~1 .lut_mask = 16'h88A8;
defparam \care_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N28
cycloneive_lcell_comb \care_ID~2 (
// Equation(s):
// \care_ID~2_combout  = (!\branch~0_combout  & \care_ID~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(\care_ID~1_combout ),
	.cin(gnd),
	.combout(\care_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \care_ID~2 .lut_mask = 16'h0F00;
defparam \care_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N2
cycloneive_lcell_comb \ALUOP_ID~0 (
// Equation(s):
// \ALUOP_ID~0_combout  = (Instr_IF_4) # ((Instr_IF_3 & ((!WideOr41))) # (!Instr_IF_3 & (WideOr4)))

	.dataa(WideOr4),
	.datab(WideOr41),
	.datac(Instr_IF_4),
	.datad(Instr_IF_3),
	.cin(gnd),
	.combout(\ALUOP_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~0 .lut_mask = 16'hF3FA;
defparam \ALUOP_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N28
cycloneive_lcell_comb \ALUOP_ID~1 (
// Equation(s):
// \ALUOP_ID~1_combout  = (Instr_IF_28 & (!Instr_IF_26 & ((Instr_IF_27)))) # (!Instr_IF_28 & (Instr_IF_26 & (Instr_IF_31)))

	.dataa(Instr_IF_28),
	.datab(Instr_IF_26),
	.datac(Instr_IF_31),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(\ALUOP_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~1 .lut_mask = 16'h6240;
defparam \ALUOP_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N20
cycloneive_lcell_comb \ALUOP_ID~2 (
// Equation(s):
// \ALUOP_ID~2_combout  = (!Instr_IF_30 & ((\ALUOP_ID~1_combout ) # (Instr_IF_28 $ (Instr_IF_29))))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_28),
	.datac(Instr_IF_29),
	.datad(\ALUOP_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUOP_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~2 .lut_mask = 16'h5514;
defparam \ALUOP_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N24
cycloneive_lcell_comb \ALUOP_ID~3 (
// Equation(s):
// \ALUOP_ID~3_combout  = (!\branch~0_combout  & ((Selector11 & ((\ALUOP_ID~2_combout ))) # (!Selector11 & (\ALUOP_ID~0_combout ))))

	.dataa(\ALUOP_ID~0_combout ),
	.datab(Selector111),
	.datac(\ALUOP_ID~2_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUOP_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~3 .lut_mask = 16'h00E2;
defparam \ALUOP_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N8
cycloneive_lcell_comb \ALUOP_ID~4 (
// Equation(s):
// \ALUOP_ID~4_combout  = (!Instr_IF_3 & (!Instr_IF_5 & ((Instr_IF_0) # (Instr_IF_2))))

	.dataa(Instr_IF_3),
	.datab(Instr_IF_5),
	.datac(Instr_IF_0),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(\ALUOP_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~4 .lut_mask = 16'h1110;
defparam \ALUOP_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N6
cycloneive_lcell_comb \ALUOP_ID~5 (
// Equation(s):
// \ALUOP_ID~5_combout  = (Instr_IF_4) # ((\ALUOP_ID~4_combout ) # ((!WideOr41 & Instr_IF_3)))

	.dataa(Instr_IF_4),
	.datab(WideOr41),
	.datac(\ALUOP_ID~4_combout ),
	.datad(Instr_IF_3),
	.cin(gnd),
	.combout(\ALUOP_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~5 .lut_mask = 16'hFBFA;
defparam \ALUOP_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N18
cycloneive_lcell_comb \ALUOP_ID~6 (
// Equation(s):
// \ALUOP_ID~6_combout  = (!Instr_IF_28 & (!Instr_IF_30 & ((!Instr_IF_31) # (!Instr_IF_26))))

	.dataa(Instr_IF_28),
	.datab(Instr_IF_26),
	.datac(Instr_IF_30),
	.datad(Instr_IF_31),
	.cin(gnd),
	.combout(\ALUOP_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~6 .lut_mask = 16'h0105;
defparam \ALUOP_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N4
cycloneive_lcell_comb \ALUOP_ID~7 (
// Equation(s):
// \ALUOP_ID~7_combout  = (Instr_IF_29 & (\ALUOP_ID~6_combout  & ((Instr_IF_27)))) # (!Instr_IF_29 & (((Selector14))))

	.dataa(Instr_IF_29),
	.datab(\ALUOP_ID~6_combout ),
	.datac(Selector141),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(\ALUOP_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~7 .lut_mask = 16'hD850;
defparam \ALUOP_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N2
cycloneive_lcell_comb \ALUOP_ID~8 (
// Equation(s):
// \ALUOP_ID~8_combout  = (\ALUOP_ID~7_combout  & (!\branch~0_combout  & ((\ALUOP_ID~5_combout ) # (Instr_IF_29))))

	.dataa(\ALUOP_ID~5_combout ),
	.datab(\ALUOP_ID~7_combout ),
	.datac(branch),
	.datad(Instr_IF_29),
	.cin(gnd),
	.combout(\ALUOP_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~8 .lut_mask = 16'h0C08;
defparam \ALUOP_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N16
cycloneive_lcell_comb \ALUOP_ID~10 (
// Equation(s):
// \ALUOP_ID~10_combout  = (!Instr_IF_3 & (Instr_IF_5 & (!Instr_IF_4 & Instr_IF_2)))

	.dataa(Instr_IF_3),
	.datab(Instr_IF_5),
	.datac(Instr_IF_4),
	.datad(Instr_IF_2),
	.cin(gnd),
	.combout(\ALUOP_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~10 .lut_mask = 16'h0400;
defparam \ALUOP_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N14
cycloneive_lcell_comb \ALUOP_ID~9 (
// Equation(s):
// \ALUOP_ID~9_combout  = (!Instr_IF_30 & (Instr_IF_29 & Instr_IF_28))

	.dataa(Instr_IF_30),
	.datab(gnd),
	.datac(Instr_IF_29),
	.datad(Instr_IF_28),
	.cin(gnd),
	.combout(\ALUOP_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~9 .lut_mask = 16'h5000;
defparam \ALUOP_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N26
cycloneive_lcell_comb \ALUOP_ID~11 (
// Equation(s):
// \ALUOP_ID~11_combout  = (!\branch~0_combout  & ((\ALUOP_ID~9_combout ) # ((\ALUOP_ID~10_combout  & !Selector11))))

	.dataa(\ALUOP_ID~10_combout ),
	.datab(Selector111),
	.datac(\ALUOP_ID~9_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUOP_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~11 .lut_mask = 16'h00F2;
defparam \ALUOP_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N26
cycloneive_lcell_comb \jump_ID~5 (
// Equation(s):
// \jump_ID~5_combout  = (!Instr_IF_30 & !\branch~0_combout )

	.dataa(Instr_IF_30),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\jump_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~5 .lut_mask = 16'h0505;
defparam \jump_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N22
cycloneive_lcell_comb \RegDst_ID~2 (
// Equation(s):
// \RegDst_ID~2_combout  = (\jump_ID~5_combout  & ((Instr_IF_29 & (!Instr_IF_31)) # (!Instr_IF_29 & (Instr_IF_31 & WideOr21))))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_31),
	.datac(\jump_ID~5_combout ),
	.datad(WideOr21),
	.cin(gnd),
	.combout(\RegDst_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_ID~2 .lut_mask = 16'h6020;
defparam \RegDst_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y28_N23
dffeas \RegDst_ID[0] (
	.clk(CLK),
	.d(\RegDst_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_ID[0]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_ID[0] .is_wysiwyg = "true";
defparam \RegDst_ID[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N20
cycloneive_lcell_comb \RegDst_ID~1 (
// Equation(s):
// \RegDst_ID~1_combout  = (!Instr_IF_29 & (!Instr_IF_31 & \RegDst_ID~0_combout ))

	.dataa(gnd),
	.datab(Instr_IF_29),
	.datac(Instr_IF_31),
	.datad(\RegDst_ID~0_combout ),
	.cin(gnd),
	.combout(\RegDst_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_ID~1 .lut_mask = 16'h0300;
defparam \RegDst_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N21
dffeas \RegDst_ID[1] (
	.clk(CLK),
	.d(\RegDst_ID~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDst_ID[1]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDst_ID[1] .is_wysiwyg = "true";
defparam \RegDst_ID[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \RegDst_EX~0 (
// Equation(s):
// \RegDst_EX~0_combout  = (RegDst_ID[1]) # ((RegDst_ID[0] & ((Instr_ID_16))) # (!RegDst_ID[0] & (Instr_ID_11)))

	.dataa(Instr_ID_11),
	.datab(RegDst_ID[0]),
	.datac(Instr_ID_16),
	.datad(RegDst_ID[1]),
	.cin(gnd),
	.combout(\RegDst_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~0 .lut_mask = 16'hFFE2;
defparam \RegDst_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \RegDst_EX~1 (
// Equation(s):
// \RegDst_EX~1_combout  = (\always1~0_combout  & (\RegDst_EX~0_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(\always1~0_combout ),
	.datac(\RegDst_EX~0_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(\RegDst_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~1 .lut_mask = 16'h40C0;
defparam \RegDst_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \RegDst_EX~2 (
// Equation(s):
// \RegDst_EX~2_combout  = (RegDst_ID[1]) # ((RegDst_ID[0] & (Instr_ID_17)) # (!RegDst_ID[0] & ((Instr_ID_12))))

	.dataa(Instr_ID_17),
	.datab(RegDst_ID[1]),
	.datac(Instr_ID_12),
	.datad(RegDst_ID[0]),
	.cin(gnd),
	.combout(\RegDst_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~2 .lut_mask = 16'hEEFC;
defparam \RegDst_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \RegDst_EX~3 (
// Equation(s):
// \RegDst_EX~3_combout  = (\always1~0_combout  & (\RegDst_EX~2_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(\always1~0_combout ),
	.datad(\RegDst_EX~2_combout ),
	.cin(gnd),
	.combout(\RegDst_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~3 .lut_mask = 16'h7000;
defparam \RegDst_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \RegDst_EX~4 (
// Equation(s):
// \RegDst_EX~4_combout  = (RegDst_ID[1]) # ((RegDst_ID[0] & (Instr_ID_18)) # (!RegDst_ID[0] & ((Instr_ID_13))))

	.dataa(Instr_ID_18),
	.datab(RegDst_ID[0]),
	.datac(Instr_ID_13),
	.datad(RegDst_ID[1]),
	.cin(gnd),
	.combout(\RegDst_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~4 .lut_mask = 16'hFFB8;
defparam \RegDst_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \RegDst_EX~5 (
// Equation(s):
// \RegDst_EX~5_combout  = (\always1~0_combout  & (\RegDst_EX~4_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(\always1~0_combout ),
	.datac(\RegDst_EX~4_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(\RegDst_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~5 .lut_mask = 16'h40C0;
defparam \RegDst_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N16
cycloneive_lcell_comb \RegWen_ID~2 (
// Equation(s):
// \RegWen_ID~2_combout  = (\RegWen_ID~1_combout  & !\branch~0_combout )

	.dataa(\RegWen_ID~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegWen_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegWen_ID~2 .lut_mask = 16'h00AA;
defparam \RegWen_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y28_N17
dffeas RegWen_ID(
	.clk(CLK),
	.d(\RegWen_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\RegWen_ID~q ),
	.prn(vcc));
// synopsys translate_off
defparam RegWen_ID.is_wysiwyg = "true";
defparam RegWen_ID.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \RegWen_EX~0 (
// Equation(s):
// \RegWen_EX~0_combout  = (\always1~0_combout  & (\RegWen_ID~q  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(\always1~0_combout ),
	.datad(\RegWen_ID~q ),
	.cin(gnd),
	.combout(\RegWen_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegWen_EX~0 .lut_mask = 16'h7000;
defparam \RegWen_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \RegDst_EX~6 (
// Equation(s):
// \RegDst_EX~6_combout  = (RegDst_ID[1]) # ((RegDst_ID[0] & (Instr_ID_19)) # (!RegDst_ID[0] & ((Instr_ID_14))))

	.dataa(Instr_ID_19),
	.datab(RegDst_ID[1]),
	.datac(RegDst_ID[0]),
	.datad(Instr_ID_14),
	.cin(gnd),
	.combout(\RegDst_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~6 .lut_mask = 16'hEFEC;
defparam \RegDst_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \RegDst_EX~7 (
// Equation(s):
// \RegDst_EX~7_combout  = (\always1~0_combout  & (\RegDst_EX~6_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(\always1~0_combout ),
	.datac(\RegDst_EX~6_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(\RegDst_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~7 .lut_mask = 16'h40C0;
defparam \RegDst_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \RegDst_EX~8 (
// Equation(s):
// \RegDst_EX~8_combout  = (RegDst_ID[1]) # ((RegDst_ID[0] & (Instr_ID_20)) # (!RegDst_ID[0] & ((Instr_ID_15))))

	.dataa(Instr_ID_20),
	.datab(RegDst_ID[0]),
	.datac(Instr_ID_15),
	.datad(RegDst_ID[1]),
	.cin(gnd),
	.combout(\RegDst_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~8 .lut_mask = 16'hFFB8;
defparam \RegDst_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \RegDst_EX~9 (
// Equation(s):
// \RegDst_EX~9_combout  = (\always1~0_combout  & (\RegDst_EX~8_combout  & ((!always01) # (!src2_hazard_t1))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(\always1~0_combout ),
	.datad(\RegDst_EX~8_combout ),
	.cin(gnd),
	.combout(\RegDst_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~9 .lut_mask = 16'h7000;
defparam \RegDst_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \Instr_ID~0 (
// Equation(s):
// \Instr_ID~0_combout  = (Instr_IF_16 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_16),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~0 .lut_mask = 16'h00CC;
defparam \Instr_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N18
cycloneive_lcell_comb \hazard_Reg_ID~0 (
// Equation(s):
// \hazard_Reg_ID~0_combout  = (!Instr_IF_30 & (!Instr_IF_28 & (!input_hazard_Reg_ID & !\branch~0_combout )))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_28),
	.datac(input_hazard_Reg_ID),
	.datad(branch),
	.cin(gnd),
	.combout(\hazard_Reg_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \hazard_Reg_ID~0 .lut_mask = 16'h0001;
defparam \hazard_Reg_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Instr_ID~1 (
// Equation(s):
// \Instr_ID~1_combout  = (!\branch~0_combout  & Instr_IF_17)

	.dataa(branch),
	.datab(gnd),
	.datac(gnd),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\Instr_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~1 .lut_mask = 16'h5500;
defparam \Instr_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Instr_ID~2 (
// Equation(s):
// \Instr_ID~2_combout  = (Instr_IF_18 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Instr_IF_18),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~2 .lut_mask = 16'h00F0;
defparam \Instr_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Instr_ID~3 (
// Equation(s):
// \Instr_ID~3_combout  = (Instr_IF_19 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_19),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~3 .lut_mask = 16'h00CC;
defparam \Instr_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \Memwrite_ID~0 (
// Equation(s):
// \Memwrite_ID~0_combout  = (Instr_IF_31 & (Instr_IF_29 & \RegDst_ID~0_combout ))

	.dataa(Instr_IF_31),
	.datab(Instr_IF_29),
	.datac(gnd),
	.datad(\RegDst_ID~0_combout ),
	.cin(gnd),
	.combout(\Memwrite_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \Memwrite_ID~0 .lut_mask = 16'h8800;
defparam \Memwrite_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \Instr_ID~4 (
// Equation(s):
// \Instr_ID~4_combout  = (!\branch~0_combout  & Instr_IF_20)

	.dataa(branch),
	.datab(gnd),
	.datac(Instr_IF_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~4 .lut_mask = 16'h5050;
defparam \Instr_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \MemToReg_MEM~feeder (
// Equation(s):
// \MemToReg_MEM~feeder_combout  = MemToReg_EX1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(MemToReg_EX1),
	.cin(gnd),
	.combout(\MemToReg_MEM~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \MemToReg_MEM~feeder .lut_mask = 16'hFF00;
defparam \MemToReg_MEM~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = (!\Equal20~0_combout  & (src2_hazard_t2 & (!src2_hazard_t1 & !always01)))

	.dataa(Equal20),
	.datab(src2_hazard_t1),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0004;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \ALUSrc2_ID~1 (
// Equation(s):
// \ALUSrc2_ID~1_combout  = (WideOr212 & (Instr_IF[15])) # (!WideOr212 & (((!WideOr14 & rfifrdat2_31))))

	.dataa(Instr_IF[15]),
	.datab(WideOr14),
	.datac(rfifrdat2_31),
	.datad(WideOr212),
	.cin(gnd),
	.combout(\ALUSrc2_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~1 .lut_mask = 16'hAA30;
defparam \ALUSrc2_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \ALUSrc2_ID~0 (
// Equation(s):
// \ALUSrc2_ID~0_combout  = (!Selector141 & (!\Equal3~0_combout  & !\branch~0_combout ))

	.dataa(Selector142),
	.datab(gnd),
	.datac(\Equal3~0_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~0 .lut_mask = 16'h0005;
defparam \ALUSrc2_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \ALUSrc2_ID~2 (
// Equation(s):
// \ALUSrc2_ID~2_combout  = (\Equal3~0_combout  & ((ReadData_MEM_31) # ((\ALUSrc2_ID~1_combout  & \ALUSrc2_ID~0_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~1_combout  & \ALUSrc2_ID~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_31),
	.datac(\ALUSrc2_ID~1_combout ),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~2 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \ALUSrc2_ID[31]~3 (
// Equation(s):
// \ALUSrc2_ID[31]~3_combout  = (always1 & ((\Equal3~0_combout ) # (!\always1~2_combout )))

	.dataa(\Equal3~0_combout ),
	.datab(\always1~2_combout ),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc2_ID[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID[31]~3 .lut_mask = 16'hB0B0;
defparam \ALUSrc2_ID[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \Instr_ID~5 (
// Equation(s):
// \Instr_ID~5_combout  = (Instr_IF_21 & !\branch~0_combout )

	.dataa(Instr_IF_21),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~5 .lut_mask = 16'h0A0A;
defparam \Instr_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Instr_ID~6 (
// Equation(s):
// \Instr_ID~6_combout  = (Instr_IF_22 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_22),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~6 .lut_mask = 16'h00CC;
defparam \Instr_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Instr_ID~7 (
// Equation(s):
// \Instr_ID~7_combout  = (Instr_IF_24 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_24),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~7 .lut_mask = 16'h00CC;
defparam \Instr_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \Instr_ID~8 (
// Equation(s):
// \Instr_ID~8_combout  = (!\branch~0_combout  & Instr_IF_25)

	.dataa(gnd),
	.datab(branch),
	.datac(gnd),
	.datad(Instr_IF_25),
	.cin(gnd),
	.combout(\Instr_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~8 .lut_mask = 16'h3300;
defparam \Instr_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Instr_ID~9 (
// Equation(s):
// \Instr_ID~9_combout  = (Instr_IF_23 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Instr_IF_23),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~9 .lut_mask = 16'h00F0;
defparam \Instr_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \ALUSrc1_ID~0 (
// Equation(s):
// \ALUSrc1_ID~0_combout  = (Instr_IF_25 & ((rfifrdat1_31))) # (!Instr_IF_25 & (rfifrdat1_311))

	.dataa(gnd),
	.datab(rfifrdat1_311),
	.datac(Instr_IF_25),
	.datad(rfifrdat1_31),
	.cin(gnd),
	.combout(\ALUSrc1_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~0 .lut_mask = 16'hFC0C;
defparam \ALUSrc1_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \ALUSrc1_ID~1 (
// Equation(s):
// \ALUSrc1_ID~1_combout  = (!\Equal20~0_combout  & (!\branch~0_combout  & ((Instr_IF_21) # (WideOr0))))

	.dataa(Instr_IF_21),
	.datab(WideOr0),
	.datac(Equal20),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc1_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~1 .lut_mask = 16'h000E;
defparam \ALUSrc1_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \ALUSrc1_ID~2 (
// Equation(s):
// \ALUSrc1_ID~2_combout  = (ReadData_MEM_31 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~0_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_31 & (\ALUSrc1_ID~0_combout  & (\ALUSrc1_ID~1_combout )))

	.dataa(ReadData_MEM_31),
	.datab(\ALUSrc1_ID~0_combout ),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(Equal20),
	.cin(gnd),
	.combout(\ALUSrc1_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~2 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \ALUSrc1_ID[31]~3 (
// Equation(s):
// \ALUSrc1_ID[31]~3_combout  = (always1 & ((\Equal20~0_combout ) # (!\always1~2_combout )))

	.dataa(always1),
	.datab(gnd),
	.datac(Equal20),
	.datad(\always1~2_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID[31]~3 .lut_mask = 16'hA0AA;
defparam \ALUSrc1_ID[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N4
cycloneive_lcell_comb \ALUOP_ID~14 (
// Equation(s):
// \ALUOP_ID~14_combout  = (Instr_IF_4) # ((Instr_IF_0 & (!WideOr61)) # (!Instr_IF_0 & ((WideOr6))))

	.dataa(Instr_IF_0),
	.datab(Instr_IF_4),
	.datac(WideOr61),
	.datad(WideOr6),
	.cin(gnd),
	.combout(\ALUOP_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~14 .lut_mask = 16'hDFCE;
defparam \ALUOP_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N16
cycloneive_lcell_comb \ALUOP_ID~12 (
// Equation(s):
// \ALUOP_ID~12_combout  = (Instr_IF_29 & (Instr_IF_26 & (!Instr_IF_31 & Instr_IF_27)))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_26),
	.datac(Instr_IF_31),
	.datad(Instr_IF_27),
	.cin(gnd),
	.combout(\ALUOP_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~12 .lut_mask = 16'h0800;
defparam \ALUOP_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N6
cycloneive_lcell_comb \ALUOP_ID~13 (
// Equation(s):
// \ALUOP_ID~13_combout  = (\ALUOP_ID~12_combout ) # ((Instr_IF_28 & ((Instr_IF_26) # (!Instr_IF_29))))

	.dataa(Instr_IF_29),
	.datab(Instr_IF_26),
	.datac(Instr_IF_28),
	.datad(\ALUOP_ID~12_combout ),
	.cin(gnd),
	.combout(\ALUOP_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~13 .lut_mask = 16'hFFD0;
defparam \ALUOP_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N12
cycloneive_lcell_comb \ALUOP_ID~15 (
// Equation(s):
// \ALUOP_ID~15_combout  = (Instr_IF_30 & (!Selector11 & (\ALUOP_ID~14_combout ))) # (!Instr_IF_30 & ((\ALUOP_ID~13_combout ) # ((!Selector11 & \ALUOP_ID~14_combout ))))

	.dataa(Instr_IF_30),
	.datab(Selector111),
	.datac(\ALUOP_ID~14_combout ),
	.datad(\ALUOP_ID~13_combout ),
	.cin(gnd),
	.combout(\ALUOP_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~15 .lut_mask = 16'h7530;
defparam \ALUOP_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N6
cycloneive_lcell_comb \ALUOP_ID~16 (
// Equation(s):
// \ALUOP_ID~16_combout  = (!\branch~0_combout  & \ALUOP_ID~15_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(\ALUOP_ID~15_combout ),
	.cin(gnd),
	.combout(\ALUOP_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ID~16 .lut_mask = 16'h0F00;
defparam \ALUOP_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \ALUSrc1_ID~4 (
// Equation(s):
// \ALUSrc1_ID~4_combout  = (Instr_IF_25 & (rfifrdat1_30)) # (!Instr_IF_25 & ((rfifrdat1_301)))

	.dataa(rfifrdat1_30),
	.datab(Instr_IF_25),
	.datac(gnd),
	.datad(rfifrdat1_301),
	.cin(gnd),
	.combout(\ALUSrc1_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~4 .lut_mask = 16'hBB88;
defparam \ALUSrc1_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \ALUSrc1_ID~5 (
// Equation(s):
// \ALUSrc1_ID~5_combout  = (\Equal20~0_combout  & ((ReadData_MEM_30) # ((\ALUSrc1_ID~4_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~4_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_30),
	.datac(\ALUSrc1_ID~4_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~5 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \ReadData_MEM[30]~feeder (
// Equation(s):
// \ReadData_MEM[30]~feeder_combout  = ramiframload_30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\ReadData_MEM[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[30]~feeder .lut_mask = 16'hFF00;
defparam \ReadData_MEM[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \Instr_IF~17 (
// Equation(s):
// \Instr_IF~17_combout  = (always1 & (!always0 & (ramiframload_15 & !\branch~0_combout )))

	.dataa(always1),
	.datab(always02),
	.datac(ramiframload_15),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~17_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~17 .lut_mask = 16'h0020;
defparam \Instr_IF~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N21
dffeas \Instr_IF[15] (
	.clk(CLK),
	.d(\Instr_IF~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF[15]),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[15] .is_wysiwyg = "true";
defparam \Instr_IF[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \ALUSrc2_ID~4 (
// Equation(s):
// \ALUSrc2_ID~4_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_30)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_30),
	.cin(gnd),
	.combout(\ALUSrc2_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~4 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \ALUSrc2_ID~5 (
// Equation(s):
// \ALUSrc2_ID~5_combout  = (\ALUSrc2_ID~4_combout ) # ((Instr_IF[14] & (WideOr212 & WideOr14)))

	.dataa(Instr_IF[14]),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(\ALUSrc2_ID~4_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~5 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \ALUSrc2_ID~6 (
// Equation(s):
// \ALUSrc2_ID~6_combout  = (ReadData_MEM_30 & ((\Equal3~0_combout ) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~5_combout )))) # (!ReadData_MEM_30 & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~5_combout ))))

	.dataa(ReadData_MEM_30),
	.datab(\Equal3~0_combout ),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~5_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~6 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \ALUSrc1_ID~6 (
// Equation(s):
// \ALUSrc1_ID~6_combout  = (Instr_IF_25 & ((rfifrdat1_29))) # (!Instr_IF_25 & (rfifrdat1_291))

	.dataa(Instr_IF_25),
	.datab(gnd),
	.datac(rfifrdat1_291),
	.datad(rfifrdat1_29),
	.cin(gnd),
	.combout(\ALUSrc1_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~6 .lut_mask = 16'hFA50;
defparam \ALUSrc1_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \ALUSrc1_ID~7 (
// Equation(s):
// \ALUSrc1_ID~7_combout  = (\ALUSrc1_ID~6_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_29 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~6_combout  & (ReadData_MEM_29 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~6_combout ),
	.datab(ReadData_MEM_29),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~7 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \CalcData_MEM[29]~feeder (
// Equation(s):
// \CalcData_MEM[29]~feeder_combout  = Result_EX_29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_29),
	.cin(gnd),
	.combout(\CalcData_MEM[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[29]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \Instr_IF~24 (
// Equation(s):
// \Instr_IF~24_combout  = (always1 & (!\branch~0_combout  & (!always0 & ramiframload_13)))

	.dataa(always1),
	.datab(branch),
	.datac(always02),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(\Instr_IF~24_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~24 .lut_mask = 16'h0200;
defparam \Instr_IF~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N21
dffeas \Instr_IF[13] (
	.clk(CLK),
	.d(\Instr_IF~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF[13]),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[13] .is_wysiwyg = "true";
defparam \Instr_IF[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \ALUSrc2_ID~7 (
// Equation(s):
// \ALUSrc2_ID~7_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_29)))))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF[15]),
	.datad(rfifrdat2_29),
	.cin(gnd),
	.combout(\ALUSrc2_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~7 .lut_mask = 16'h5140;
defparam \ALUSrc2_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \ALUSrc2_ID~8 (
// Equation(s):
// \ALUSrc2_ID~8_combout  = (\ALUSrc2_ID~7_combout ) # ((WideOr14 & (WideOr212 & Instr_IF[13])))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF[13]),
	.datad(\ALUSrc2_ID~7_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~8 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \ALUSrc2_ID~9 (
// Equation(s):
// \ALUSrc2_ID~9_combout  = (\ALUSrc2_ID~8_combout  & ((\ALUSrc2_ID~0_combout ) # ((ReadData_MEM_29 & \Equal3~0_combout )))) # (!\ALUSrc2_ID~8_combout  & (ReadData_MEM_29 & (\Equal3~0_combout )))

	.dataa(\ALUSrc2_ID~8_combout ),
	.datab(ReadData_MEM_29),
	.datac(\Equal3~0_combout ),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~9 .lut_mask = 16'hEAC0;
defparam \ALUSrc2_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \ALUSrc1_ID~8 (
// Equation(s):
// \ALUSrc1_ID~8_combout  = (Instr_IF_25 & ((rfifrdat1_28))) # (!Instr_IF_25 & (rfifrdat1_281))

	.dataa(rfifrdat1_281),
	.datab(Instr_IF_25),
	.datac(gnd),
	.datad(rfifrdat1_28),
	.cin(gnd),
	.combout(\ALUSrc1_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~8 .lut_mask = 16'hEE22;
defparam \ALUSrc1_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \ALUSrc1_ID~9 (
// Equation(s):
// \ALUSrc1_ID~9_combout  = (\Equal20~0_combout  & ((ReadData_MEM_28) # ((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~8_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~8_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_28),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(\ALUSrc1_ID~8_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~9 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N28
cycloneive_lcell_comb \Instr_IF~25 (
// Equation(s):
// \Instr_IF~25_combout  = (!always0 & (!\branch~0_combout  & (always1 & ramiframload_12)))

	.dataa(always02),
	.datab(branch),
	.datac(always1),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(\Instr_IF~25_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~25 .lut_mask = 16'h1000;
defparam \Instr_IF~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N29
dffeas \Instr_IF[12] (
	.clk(CLK),
	.d(\Instr_IF~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF[12]),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[12] .is_wysiwyg = "true";
defparam \Instr_IF[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \ALUSrc2_ID~10 (
// Equation(s):
// \ALUSrc2_ID~10_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_28)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_28),
	.cin(gnd),
	.combout(\ALUSrc2_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~10 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \ALUSrc2_ID~11 (
// Equation(s):
// \ALUSrc2_ID~11_combout  = (\ALUSrc2_ID~10_combout ) # ((WideOr14 & (WideOr212 & Instr_IF[12])))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF[12]),
	.datad(\ALUSrc2_ID~10_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~11 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \ALUSrc2_ID~12 (
// Equation(s):
// \ALUSrc2_ID~12_combout  = (ReadData_MEM_28 & ((\Equal3~0_combout ) # ((\ALUSrc2_ID~11_combout  & \ALUSrc2_ID~0_combout )))) # (!ReadData_MEM_28 & (((\ALUSrc2_ID~11_combout  & \ALUSrc2_ID~0_combout ))))

	.dataa(ReadData_MEM_28),
	.datab(\Equal3~0_combout ),
	.datac(\ALUSrc2_ID~11_combout ),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~12 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \ALUSrc1_ID~10 (
// Equation(s):
// \ALUSrc1_ID~10_combout  = (Instr_IF_25 & ((rfifrdat1_27))) # (!Instr_IF_25 & (rfifrdat1_271))

	.dataa(rfifrdat1_271),
	.datab(rfifrdat1_27),
	.datac(gnd),
	.datad(Instr_IF_25),
	.cin(gnd),
	.combout(\ALUSrc1_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~10 .lut_mask = 16'hCCAA;
defparam \ALUSrc1_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \ALUSrc1_ID~11 (
// Equation(s):
// \ALUSrc1_ID~11_combout  = (\ALUSrc1_ID~10_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_27 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~10_combout  & (ReadData_MEM_27 & ((\Equal20~0_combout ))))

	.dataa(\ALUSrc1_ID~10_combout ),
	.datab(ReadData_MEM_27),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(Equal20),
	.cin(gnd),
	.combout(\ALUSrc1_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~11 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \ReadData_MEM[27]~feeder (
// Equation(s):
// \ReadData_MEM[27]~feeder_combout  = ramiframload_27

	.dataa(gnd),
	.datab(ramiframload_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[27]~feeder .lut_mask = 16'hCCCC;
defparam \ReadData_MEM[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N16
cycloneive_lcell_comb \Instr_IF~26 (
// Equation(s):
// \Instr_IF~26_combout  = (ramiframload_11 & (!always0 & (!\branch~0_combout  & always1)))

	.dataa(ramiframload_11),
	.datab(always02),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~26_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~26 .lut_mask = 16'h0200;
defparam \Instr_IF~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N17
dffeas \Instr_IF[11] (
	.clk(CLK),
	.d(\Instr_IF~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF[11]),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[11] .is_wysiwyg = "true";
defparam \Instr_IF[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N2
cycloneive_lcell_comb \ALUSrc2_ID~13 (
// Equation(s):
// \ALUSrc2_ID~13_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_27)))))

	.dataa(Instr_IF[15]),
	.datab(WideOr14),
	.datac(rfifrdat2_27),
	.datad(WideOr212),
	.cin(gnd),
	.combout(\ALUSrc2_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~13 .lut_mask = 16'h2230;
defparam \ALUSrc2_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \ALUSrc2_ID~14 (
// Equation(s):
// \ALUSrc2_ID~14_combout  = (\ALUSrc2_ID~13_combout ) # ((WideOr212 & (WideOr14 & Instr_IF[11])))

	.dataa(WideOr212),
	.datab(WideOr14),
	.datac(Instr_IF[11]),
	.datad(\ALUSrc2_ID~13_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~14 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \ALUSrc2_ID~15 (
// Equation(s):
// \ALUSrc2_ID~15_combout  = (\Equal3~0_combout  & ((ReadData_MEM_27) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~14_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~14_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_27),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~14_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~15 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \ALUSrc1_ID~12 (
// Equation(s):
// \ALUSrc1_ID~12_combout  = (Instr_IF_25 & ((rfifrdat1_26))) # (!Instr_IF_25 & (rfifrdat1_261))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_261),
	.datac(gnd),
	.datad(rfifrdat1_26),
	.cin(gnd),
	.combout(\ALUSrc1_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~12 .lut_mask = 16'hEE44;
defparam \ALUSrc1_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \ALUSrc1_ID~13 (
// Equation(s):
// \ALUSrc1_ID~13_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~12_combout ) # ((ReadData_MEM_26 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~1_combout  & (ReadData_MEM_26 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(ReadData_MEM_26),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~12_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~13 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \CalcData_MEM[26]~feeder (
// Equation(s):
// \CalcData_MEM[26]~feeder_combout  = Result_EX_26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_26),
	.cin(gnd),
	.combout(\CalcData_MEM[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[26]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \ALUSrc2_ID~16 (
// Equation(s):
// \ALUSrc2_ID~16_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_26)))))

	.dataa(Instr_IF[15]),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(rfifrdat2_26),
	.cin(gnd),
	.combout(\ALUSrc2_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~16 .lut_mask = 16'h0B08;
defparam \ALUSrc2_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \ALUSrc2_ID~17 (
// Equation(s):
// \ALUSrc2_ID~17_combout  = (\ALUSrc2_ID~16_combout ) # ((Instr_IF_10 & (WideOr212 & WideOr14)))

	.dataa(Instr_IF_10),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(\ALUSrc2_ID~16_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~17_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~17 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N14
cycloneive_lcell_comb \ALUSrc2_ID~18 (
// Equation(s):
// \ALUSrc2_ID~18_combout  = (\Equal3~0_combout  & ((ReadData_MEM_26) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~17_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~17_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_26),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~17_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~18_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~18 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \ALUSrc1_ID~14 (
// Equation(s):
// \ALUSrc1_ID~14_combout  = (Instr_IF_25 & (rfifrdat1_25)) # (!Instr_IF_25 & ((rfifrdat1_251)))

	.dataa(rfifrdat1_25),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_251),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc1_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~14 .lut_mask = 16'hB8B8;
defparam \ALUSrc1_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \ALUSrc1_ID~15 (
// Equation(s):
// \ALUSrc1_ID~15_combout  = (\ALUSrc1_ID~14_combout  & ((\ALUSrc1_ID~1_combout ) # ((\Equal20~0_combout  & ReadData_MEM_25)))) # (!\ALUSrc1_ID~14_combout  & (\Equal20~0_combout  & (ReadData_MEM_25)))

	.dataa(\ALUSrc1_ID~14_combout ),
	.datab(Equal20),
	.datac(ReadData_MEM_25),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~15 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N26
cycloneive_lcell_comb \ReadData_MEM[25]~feeder (
// Equation(s):
// \ReadData_MEM[25]~feeder_combout  = ramiframload_25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(\ReadData_MEM[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[25]~feeder .lut_mask = 16'hFF00;
defparam \ReadData_MEM[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \ALUSrc2_ID~19 (
// Equation(s):
// \ALUSrc2_ID~19_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_25)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_25),
	.cin(gnd),
	.combout(\ALUSrc2_ID~19_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~19 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \ALUSrc2_ID~20 (
// Equation(s):
// \ALUSrc2_ID~20_combout  = (\ALUSrc2_ID~19_combout ) # ((WideOr212 & (Instr_IF_9 & WideOr14)))

	.dataa(WideOr212),
	.datab(\ALUSrc2_ID~19_combout ),
	.datac(Instr_IF_9),
	.datad(WideOr14),
	.cin(gnd),
	.combout(\ALUSrc2_ID~20_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~20 .lut_mask = 16'hECCC;
defparam \ALUSrc2_ID~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \ALUSrc2_ID~21 (
// Equation(s):
// \ALUSrc2_ID~21_combout  = (\Equal3~0_combout  & ((ReadData_MEM_25) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~20_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~20_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_25),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~20_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~21_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~21 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \ALUSrc1_ID~16 (
// Equation(s):
// \ALUSrc1_ID~16_combout  = (Instr_IF_25 & ((rfifrdat1_24))) # (!Instr_IF_25 & (rfifrdat1_241))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_241),
	.datac(gnd),
	.datad(rfifrdat1_24),
	.cin(gnd),
	.combout(\ALUSrc1_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~16 .lut_mask = 16'hEE44;
defparam \ALUSrc1_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \ALUSrc1_ID~17 (
// Equation(s):
// \ALUSrc1_ID~17_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~16_combout ) # ((\Equal20~0_combout  & ReadData_MEM_24)))) # (!\ALUSrc1_ID~1_combout  & (\Equal20~0_combout  & (ReadData_MEM_24)))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(Equal20),
	.datac(ReadData_MEM_24),
	.datad(\ALUSrc1_ID~16_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~17_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~17 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \ALUSrc2_ID~22 (
// Equation(s):
// \ALUSrc2_ID~22_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_24)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_24),
	.cin(gnd),
	.combout(\ALUSrc2_ID~22_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~22 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \ALUSrc2_ID~23 (
// Equation(s):
// \ALUSrc2_ID~23_combout  = (\ALUSrc2_ID~22_combout ) # ((Instr_IF_8 & (WideOr212 & WideOr14)))

	.dataa(Instr_IF_8),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(\ALUSrc2_ID~22_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~23_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~23 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \ALUSrc2_ID~24 (
// Equation(s):
// \ALUSrc2_ID~24_combout  = (\Equal3~0_combout  & ((ReadData_MEM_24) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~23_combout )))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~0_combout  & ((\ALUSrc2_ID~23_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(\ALUSrc2_ID~0_combout ),
	.datac(ReadData_MEM_24),
	.datad(\ALUSrc2_ID~23_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~24_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~24 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \ALUSrc1_ID~18 (
// Equation(s):
// \ALUSrc1_ID~18_combout  = (Instr_IF_25 & (rfifrdat1_23)) # (!Instr_IF_25 & ((rfifrdat1_231)))

	.dataa(rfifrdat1_23),
	.datab(Instr_IF_25),
	.datac(gnd),
	.datad(rfifrdat1_231),
	.cin(gnd),
	.combout(\ALUSrc1_ID~18_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~18 .lut_mask = 16'hBB88;
defparam \ALUSrc1_ID~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \ALUSrc1_ID~19 (
// Equation(s):
// \ALUSrc1_ID~19_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~18_combout ) # ((ReadData_MEM_23 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~1_combout  & (ReadData_MEM_23 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(ReadData_MEM_23),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~18_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~19_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~19 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \ALUSrc2_ID~25 (
// Equation(s):
// \ALUSrc2_ID~25_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_23)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_23),
	.cin(gnd),
	.combout(\ALUSrc2_ID~25_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~25 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \ALUSrc2_ID~26 (
// Equation(s):
// \ALUSrc2_ID~26_combout  = (\ALUSrc2_ID~25_combout ) # ((WideOr212 & (WideOr14 & Instr_IF_7)))

	.dataa(WideOr212),
	.datab(WideOr14),
	.datac(\ALUSrc2_ID~25_combout ),
	.datad(Instr_IF_7),
	.cin(gnd),
	.combout(\ALUSrc2_ID~26_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~26 .lut_mask = 16'hF8F0;
defparam \ALUSrc2_ID~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \ALUSrc2_ID~27 (
// Equation(s):
// \ALUSrc2_ID~27_combout  = (ReadData_MEM_23 & ((\Equal3~0_combout ) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~26_combout )))) # (!ReadData_MEM_23 & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~26_combout ))))

	.dataa(ReadData_MEM_23),
	.datab(\Equal3~0_combout ),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~26_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~27_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~27 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \ALUSrc1_ID~20 (
// Equation(s):
// \ALUSrc1_ID~20_combout  = (Instr_IF_25 & ((rfifrdat1_22))) # (!Instr_IF_25 & (rfifrdat1_221))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_221),
	.datac(rfifrdat1_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc1_ID~20_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~20 .lut_mask = 16'hE4E4;
defparam \ALUSrc1_ID~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \ALUSrc1_ID~21 (
// Equation(s):
// \ALUSrc1_ID~21_combout  = (\ALUSrc1_ID~20_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_22 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~20_combout  & (ReadData_MEM_22 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~20_combout ),
	.datab(ReadData_MEM_22),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~21_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~21 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \ReadData_MEM[22]~feeder (
// Equation(s):
// \ReadData_MEM[22]~feeder_combout  = ramiframload_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\ReadData_MEM[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[22]~feeder .lut_mask = 16'hFF00;
defparam \ReadData_MEM[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \CalcData_MEM[22]~feeder (
// Equation(s):
// \CalcData_MEM[22]~feeder_combout  = Result_EX_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_22),
	.cin(gnd),
	.combout(\CalcData_MEM[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[22]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \ALUSrc2_ID~28 (
// Equation(s):
// \ALUSrc2_ID~28_combout  = (!WideOr14 & ((WideOr212 & ((Instr_IF[15]))) # (!WideOr212 & (rfifrdat2_22))))

	.dataa(WideOr212),
	.datab(WideOr14),
	.datac(rfifrdat2_22),
	.datad(Instr_IF[15]),
	.cin(gnd),
	.combout(\ALUSrc2_ID~28_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~28 .lut_mask = 16'h3210;
defparam \ALUSrc2_ID~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \ALUSrc2_ID~29 (
// Equation(s):
// \ALUSrc2_ID~29_combout  = (\ALUSrc2_ID~28_combout ) # ((WideOr212 & (WideOr14 & Instr_IF_6)))

	.dataa(WideOr212),
	.datab(WideOr14),
	.datac(\ALUSrc2_ID~28_combout ),
	.datad(Instr_IF_6),
	.cin(gnd),
	.combout(\ALUSrc2_ID~29_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~29 .lut_mask = 16'hF8F0;
defparam \ALUSrc2_ID~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \ALUSrc2_ID~30 (
// Equation(s):
// \ALUSrc2_ID~30_combout  = (\Equal3~0_combout  & ((ReadData_MEM_22) # ((\ALUSrc2_ID~29_combout  & \ALUSrc2_ID~0_combout )))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~29_combout  & ((\ALUSrc2_ID~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(\ALUSrc2_ID~29_combout ),
	.datac(ReadData_MEM_22),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~30_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~30 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \ALUSrc1_ID~22 (
// Equation(s):
// \ALUSrc1_ID~22_combout  = (Instr_IF_25 & ((rfifrdat1_21))) # (!Instr_IF_25 & (rfifrdat1_211))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_211),
	.datad(rfifrdat1_21),
	.cin(gnd),
	.combout(\ALUSrc1_ID~22_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~22 .lut_mask = 16'hFC30;
defparam \ALUSrc1_ID~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \ALUSrc1_ID~23 (
// Equation(s):
// \ALUSrc1_ID~23_combout  = (ReadData_MEM_21 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~22_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_21 & (\ALUSrc1_ID~22_combout  & ((\ALUSrc1_ID~1_combout ))))

	.dataa(ReadData_MEM_21),
	.datab(\ALUSrc1_ID~22_combout ),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~23_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~23 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \ReadData_MEM[21]~feeder (
// Equation(s):
// \ReadData_MEM[21]~feeder_combout  = ramiframload_21

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[21]~feeder .lut_mask = 16'hF0F0;
defparam \ReadData_MEM[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \CalcData_MEM[21]~feeder (
// Equation(s):
// \CalcData_MEM[21]~feeder_combout  = Result_EX_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_21),
	.cin(gnd),
	.combout(\CalcData_MEM[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[21]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \ALUSrc2_ID~31 (
// Equation(s):
// \ALUSrc2_ID~31_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_21)))))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF[15]),
	.datad(rfifrdat2_21),
	.cin(gnd),
	.combout(\ALUSrc2_ID~31_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~31 .lut_mask = 16'h5140;
defparam \ALUSrc2_ID~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \ALUSrc2_ID~32 (
// Equation(s):
// \ALUSrc2_ID~32_combout  = (\ALUSrc2_ID~31_combout ) # ((Instr_IF_5 & (WideOr212 & WideOr14)))

	.dataa(Instr_IF_5),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(\ALUSrc2_ID~31_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~32_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~32 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \ALUSrc2_ID~33 (
// Equation(s):
// \ALUSrc2_ID~33_combout  = (ReadData_MEM_21 & ((\Equal3~0_combout ) # ((\ALUSrc2_ID~32_combout  & \ALUSrc2_ID~0_combout )))) # (!ReadData_MEM_21 & (\ALUSrc2_ID~32_combout  & ((\ALUSrc2_ID~0_combout ))))

	.dataa(ReadData_MEM_21),
	.datab(\ALUSrc2_ID~32_combout ),
	.datac(\Equal3~0_combout ),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~33_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~33 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \ALUSrc1_ID~24 (
// Equation(s):
// \ALUSrc1_ID~24_combout  = (Instr_IF_25 & (rfifrdat1_20)) # (!Instr_IF_25 & ((rfifrdat1_201)))

	.dataa(rfifrdat1_20),
	.datab(rfifrdat1_201),
	.datac(gnd),
	.datad(Instr_IF_25),
	.cin(gnd),
	.combout(\ALUSrc1_ID~24_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~24 .lut_mask = 16'hAACC;
defparam \ALUSrc1_ID~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \ALUSrc1_ID~25 (
// Equation(s):
// \ALUSrc1_ID~25_combout  = (\Equal20~0_combout  & ((ReadData_MEM_20) # ((\ALUSrc1_ID~24_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~24_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_20),
	.datac(\ALUSrc1_ID~24_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~25_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~25 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \ReadData_MEM[20]~feeder (
// Equation(s):
// \ReadData_MEM[20]~feeder_combout  = ramiframload_20

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[20]~feeder .lut_mask = 16'hF0F0;
defparam \ReadData_MEM[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \ALUSrc2_ID~34 (
// Equation(s):
// \ALUSrc2_ID~34_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_20)))))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF[15]),
	.datad(rfifrdat2_20),
	.cin(gnd),
	.combout(\ALUSrc2_ID~34_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~34 .lut_mask = 16'h5140;
defparam \ALUSrc2_ID~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \ALUSrc2_ID~35 (
// Equation(s):
// \ALUSrc2_ID~35_combout  = (\ALUSrc2_ID~34_combout ) # ((WideOr14 & (WideOr212 & Instr_IF_4)))

	.dataa(WideOr14),
	.datab(WideOr212),
	.datac(Instr_IF_4),
	.datad(\ALUSrc2_ID~34_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~35_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~35 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \ALUSrc2_ID~36 (
// Equation(s):
// \ALUSrc2_ID~36_combout  = (ReadData_MEM_20 & ((\Equal3~0_combout ) # ((\ALUSrc2_ID~35_combout  & \ALUSrc2_ID~0_combout )))) # (!ReadData_MEM_20 & (\ALUSrc2_ID~35_combout  & ((\ALUSrc2_ID~0_combout ))))

	.dataa(ReadData_MEM_20),
	.datab(\ALUSrc2_ID~35_combout ),
	.datac(\Equal3~0_combout ),
	.datad(\ALUSrc2_ID~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~36_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~36 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \ALUSrc1_ID~26 (
// Equation(s):
// \ALUSrc1_ID~26_combout  = (Instr_IF_25 & ((rfifrdat1_19))) # (!Instr_IF_25 & (rfifrdat1_191))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_191),
	.datad(rfifrdat1_19),
	.cin(gnd),
	.combout(\ALUSrc1_ID~26_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~26 .lut_mask = 16'hFC30;
defparam \ALUSrc1_ID~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \ALUSrc1_ID~27 (
// Equation(s):
// \ALUSrc1_ID~27_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~26_combout ) # ((ReadData_MEM_19 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~1_combout  & (ReadData_MEM_19 & ((\Equal20~0_combout ))))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(ReadData_MEM_19),
	.datac(\ALUSrc1_ID~26_combout ),
	.datad(Equal20),
	.cin(gnd),
	.combout(\ALUSrc1_ID~27_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~27 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \ALUSrc2_ID~37 (
// Equation(s):
// \ALUSrc2_ID~37_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_19)))))

	.dataa(Instr_IF[15]),
	.datab(rfifrdat2_19),
	.datac(WideOr212),
	.datad(WideOr14),
	.cin(gnd),
	.combout(\ALUSrc2_ID~37_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~37 .lut_mask = 16'h00AC;
defparam \ALUSrc2_ID~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \ALUSrc2_ID~38 (
// Equation(s):
// \ALUSrc2_ID~38_combout  = (\ALUSrc2_ID~37_combout ) # ((WideOr14 & (Instr_IF_3 & WideOr212)))

	.dataa(WideOr14),
	.datab(Instr_IF_3),
	.datac(WideOr212),
	.datad(\ALUSrc2_ID~37_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~38_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~38 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \ALUSrc2_ID~39 (
// Equation(s):
// \ALUSrc2_ID~39_combout  = (\ALUSrc2_ID~0_combout  & ((\ALUSrc2_ID~38_combout ) # ((\Equal3~0_combout  & ReadData_MEM_19)))) # (!\ALUSrc2_ID~0_combout  & (\Equal3~0_combout  & (ReadData_MEM_19)))

	.dataa(\ALUSrc2_ID~0_combout ),
	.datab(\Equal3~0_combout ),
	.datac(ReadData_MEM_19),
	.datad(\ALUSrc2_ID~38_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~39_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~39 .lut_mask = 16'hEAC0;
defparam \ALUSrc2_ID~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \ALUSrc1_ID~28 (
// Equation(s):
// \ALUSrc1_ID~28_combout  = (Instr_IF_25 & ((rfifrdat1_18))) # (!Instr_IF_25 & (rfifrdat1_181))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_181),
	.datad(rfifrdat1_18),
	.cin(gnd),
	.combout(\ALUSrc1_ID~28_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~28 .lut_mask = 16'hFC30;
defparam \ALUSrc1_ID~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \ALUSrc1_ID~29 (
// Equation(s):
// \ALUSrc1_ID~29_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~28_combout ) # ((\Equal20~0_combout  & ReadData_MEM_18)))) # (!\ALUSrc1_ID~1_combout  & (\Equal20~0_combout  & (ReadData_MEM_18)))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(Equal20),
	.datac(ReadData_MEM_18),
	.datad(\ALUSrc1_ID~28_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~29_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~29 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \ReadData_MEM[18]~feeder (
// Equation(s):
// \ReadData_MEM[18]~feeder_combout  = ramiframload_18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\ReadData_MEM[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[18]~feeder .lut_mask = 16'hFF00;
defparam \ReadData_MEM[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \ALUSrc2_ID~40 (
// Equation(s):
// \ALUSrc2_ID~40_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_18)))))

	.dataa(Instr_IF[15]),
	.datab(rfifrdat2_18),
	.datac(WideOr212),
	.datad(WideOr14),
	.cin(gnd),
	.combout(\ALUSrc2_ID~40_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~40 .lut_mask = 16'h00AC;
defparam \ALUSrc2_ID~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \ALUSrc2_ID~41 (
// Equation(s):
// \ALUSrc2_ID~41_combout  = (\ALUSrc2_ID~40_combout ) # ((Instr_IF_2 & (WideOr212 & WideOr14)))

	.dataa(Instr_IF_2),
	.datab(WideOr212),
	.datac(WideOr14),
	.datad(\ALUSrc2_ID~40_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~41_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~41 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \ALUSrc2_ID~42 (
// Equation(s):
// \ALUSrc2_ID~42_combout  = (\Equal3~0_combout  & ((ReadData_MEM_18) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~41_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~41_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_18),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~41_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~42_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~42 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \ALUSrc1_ID~30 (
// Equation(s):
// \ALUSrc1_ID~30_combout  = (Instr_IF_25 & ((rfifrdat1_17))) # (!Instr_IF_25 & (rfifrdat1_171))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_171),
	.datac(rfifrdat1_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc1_ID~30_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~30 .lut_mask = 16'hE4E4;
defparam \ALUSrc1_ID~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \ALUSrc1_ID~31 (
// Equation(s):
// \ALUSrc1_ID~31_combout  = (\Equal20~0_combout  & ((ReadData_MEM_17) # ((\ALUSrc1_ID~30_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~30_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_17),
	.datac(\ALUSrc1_ID~30_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~31_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~31 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \ALUSrc2_ID~43 (
// Equation(s):
// \ALUSrc2_ID~43_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_17)))))

	.dataa(WideOr14),
	.datab(Instr_IF[15]),
	.datac(WideOr212),
	.datad(rfifrdat2_17),
	.cin(gnd),
	.combout(\ALUSrc2_ID~43_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~43 .lut_mask = 16'h4540;
defparam \ALUSrc2_ID~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \ALUSrc2_ID~44 (
// Equation(s):
// \ALUSrc2_ID~44_combout  = (\ALUSrc2_ID~43_combout ) # ((WideOr14 & (Instr_IF_1 & WideOr212)))

	.dataa(WideOr14),
	.datab(Instr_IF_1),
	.datac(WideOr212),
	.datad(\ALUSrc2_ID~43_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~44_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~44 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \ALUSrc2_ID~45 (
// Equation(s):
// \ALUSrc2_ID~45_combout  = (\Equal3~0_combout  & ((ReadData_MEM_17) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~44_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~44_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_17),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~44_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~45_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~45 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \ALUSrc1_ID~32 (
// Equation(s):
// \ALUSrc1_ID~32_combout  = (Instr_IF_25 & ((rfifrdat1_16))) # (!Instr_IF_25 & (rfifrdat1_161))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_161),
	.datad(rfifrdat1_16),
	.cin(gnd),
	.combout(\ALUSrc1_ID~32_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~32 .lut_mask = 16'hFC30;
defparam \ALUSrc1_ID~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \ALUSrc1_ID~33 (
// Equation(s):
// \ALUSrc1_ID~33_combout  = (\ALUSrc1_ID~1_combout  & ((\ALUSrc1_ID~32_combout ) # ((\Equal20~0_combout  & ReadData_MEM_16)))) # (!\ALUSrc1_ID~1_combout  & (\Equal20~0_combout  & (ReadData_MEM_16)))

	.dataa(\ALUSrc1_ID~1_combout ),
	.datab(Equal20),
	.datac(ReadData_MEM_16),
	.datad(\ALUSrc1_ID~32_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~33_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~33 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \ReadData_MEM[16]~feeder (
// Equation(s):
// \ReadData_MEM[16]~feeder_combout  = ramiframload_16

	.dataa(gnd),
	.datab(ramiframload_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[16]~feeder .lut_mask = 16'hCCCC;
defparam \ReadData_MEM[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \CalcData_MEM[16]~feeder (
// Equation(s):
// \CalcData_MEM[16]~feeder_combout  = Result_EX_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_16),
	.cin(gnd),
	.combout(\CalcData_MEM[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[16]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \ALUSrc2_ID~46 (
// Equation(s):
// \ALUSrc2_ID~46_combout  = (!WideOr14 & ((WideOr212 & (Instr_IF[15])) # (!WideOr212 & ((rfifrdat2_16)))))

	.dataa(Instr_IF[15]),
	.datab(WideOr14),
	.datac(WideOr212),
	.datad(rfifrdat2_16),
	.cin(gnd),
	.combout(\ALUSrc2_ID~46_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~46 .lut_mask = 16'h2320;
defparam \ALUSrc2_ID~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \ALUSrc2_ID~47 (
// Equation(s):
// \ALUSrc2_ID~47_combout  = (\ALUSrc2_ID~46_combout ) # ((Instr_IF_0 & (WideOr14 & WideOr212)))

	.dataa(Instr_IF_0),
	.datab(WideOr14),
	.datac(WideOr212),
	.datad(\ALUSrc2_ID~46_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~47_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~47 .lut_mask = 16'hFF80;
defparam \ALUSrc2_ID~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \ALUSrc2_ID~48 (
// Equation(s):
// \ALUSrc2_ID~48_combout  = (\Equal3~0_combout  & ((ReadData_MEM_16) # ((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~47_combout )))) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~0_combout  & \ALUSrc2_ID~47_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_16),
	.datac(\ALUSrc2_ID~0_combout ),
	.datad(\ALUSrc2_ID~47_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~48_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~48 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \ALUSrc1_ID~34 (
// Equation(s):
// \ALUSrc1_ID~34_combout  = (Instr_IF_25 & ((rfifrdat1_15))) # (!Instr_IF_25 & (rfifrdat1_151))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_151),
	.datac(gnd),
	.datad(rfifrdat1_15),
	.cin(gnd),
	.combout(\ALUSrc1_ID~34_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~34 .lut_mask = 16'hEE44;
defparam \ALUSrc1_ID~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \ALUSrc1_ID~35 (
// Equation(s):
// \ALUSrc1_ID~35_combout  = (\ALUSrc1_ID~34_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_15 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~34_combout  & (ReadData_MEM_15 & ((\Equal20~0_combout ))))

	.dataa(\ALUSrc1_ID~34_combout ),
	.datab(ReadData_MEM_15),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(Equal20),
	.cin(gnd),
	.combout(\ALUSrc1_ID~35_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~35 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \CalcData_MEM[15]~feeder (
// Equation(s):
// \CalcData_MEM[15]~feeder_combout  = Result_EX_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_15),
	.cin(gnd),
	.combout(\CalcData_MEM[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[15]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \ALUSrc2_ID~49 (
// Equation(s):
// \ALUSrc2_ID~49_combout  = (!Selector141 & (WideOr14 $ (((!Instr_IF_30 & WideOr211)))))

	.dataa(Instr_IF_30),
	.datab(WideOr211),
	.datac(Selector142),
	.datad(WideOr14),
	.cin(gnd),
	.combout(\ALUSrc2_ID~49_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~49 .lut_mask = 16'h0B04;
defparam \ALUSrc2_ID~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \ALUSrc2_ID~50 (
// Equation(s):
// \ALUSrc2_ID~50_combout  = (Instr_IF[15] & ((\ALUSrc2_ID~49_combout ) # ((rfifrdat2_15 & \Equal0~0_combout )))) # (!Instr_IF[15] & (((rfifrdat2_15 & \Equal0~0_combout ))))

	.dataa(Instr_IF[15]),
	.datab(\ALUSrc2_ID~49_combout ),
	.datac(rfifrdat2_15),
	.datad(Equal0),
	.cin(gnd),
	.combout(\ALUSrc2_ID~50_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~50 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \ALUSrc2_ID~51 (
// Equation(s):
// \ALUSrc2_ID~51_combout  = (\Equal3~0_combout  & (ReadData_MEM_15)) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~50_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_15),
	.datac(\ALUSrc2_ID~50_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~51_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~51 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \ALUSrc1_ID~36 (
// Equation(s):
// \ALUSrc1_ID~36_combout  = (Instr_IF_25 & ((rfifrdat1_14))) # (!Instr_IF_25 & (rfifrdat1_141))

	.dataa(Instr_IF_25),
	.datab(gnd),
	.datac(rfifrdat1_141),
	.datad(rfifrdat1_14),
	.cin(gnd),
	.combout(\ALUSrc1_ID~36_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~36 .lut_mask = 16'hFA50;
defparam \ALUSrc1_ID~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \ALUSrc1_ID~37 (
// Equation(s):
// \ALUSrc1_ID~37_combout  = (ReadData_MEM_14 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~36_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_14 & (\ALUSrc1_ID~36_combout  & (\ALUSrc1_ID~1_combout )))

	.dataa(ReadData_MEM_14),
	.datab(\ALUSrc1_ID~36_combout ),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(Equal20),
	.cin(gnd),
	.combout(\ALUSrc1_ID~37_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~37 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N26
cycloneive_lcell_comb \ReadData_MEM[14]~feeder (
// Equation(s):
// \ReadData_MEM[14]~feeder_combout  = ramiframload_14

	.dataa(ramiframload_14),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[14]~feeder .lut_mask = 16'hAAAA;
defparam \ReadData_MEM[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \Instr_IF~23 (
// Equation(s):
// \Instr_IF~23_combout  = (ramiframload_14 & (!always0 & (!\branch~0_combout  & always1)))

	.dataa(ramiframload_14),
	.datab(always02),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~23_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~23 .lut_mask = 16'h0200;
defparam \Instr_IF~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N13
dffeas \Instr_IF[14] (
	.clk(CLK),
	.d(\Instr_IF~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(Instr_IF[14]),
	.prn(vcc));
// synopsys translate_off
defparam \Instr_IF[14] .is_wysiwyg = "true";
defparam \Instr_IF[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N18
cycloneive_lcell_comb \ALUSrc2_ID~52 (
// Equation(s):
// \ALUSrc2_ID~52_combout  = (\ALUSrc2_ID~49_combout  & ((Instr_IF[14]) # ((\Equal0~0_combout  & rfifrdat2_14)))) # (!\ALUSrc2_ID~49_combout  & (\Equal0~0_combout  & ((rfifrdat2_14))))

	.dataa(\ALUSrc2_ID~49_combout ),
	.datab(Equal0),
	.datac(Instr_IF[14]),
	.datad(rfifrdat2_14),
	.cin(gnd),
	.combout(\ALUSrc2_ID~52_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~52 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N0
cycloneive_lcell_comb \ALUSrc2_ID~53 (
// Equation(s):
// \ALUSrc2_ID~53_combout  = (\Equal3~0_combout  & (((ReadData_MEM_14)))) # (!\Equal3~0_combout  & (!\branch~0_combout  & ((\ALUSrc2_ID~52_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(branch),
	.datac(ReadData_MEM_14),
	.datad(\ALUSrc2_ID~52_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~53_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~53 .lut_mask = 16'hB1A0;
defparam \ALUSrc2_ID~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N6
cycloneive_lcell_comb \ALUSrc2_ID~54 (
// Equation(s):
// \ALUSrc2_ID~54_combout  = (Instr_IF[13] & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_13)))) # (!Instr_IF[13] & (((\Equal0~0_combout  & rfifrdat2_13))))

	.dataa(Instr_IF[13]),
	.datab(\ALUSrc2_ID~49_combout ),
	.datac(Equal0),
	.datad(rfifrdat2_13),
	.cin(gnd),
	.combout(\ALUSrc2_ID~54_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~54 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N28
cycloneive_lcell_comb \ALUSrc2_ID~55 (
// Equation(s):
// \ALUSrc2_ID~55_combout  = (\Equal3~0_combout  & (ReadData_MEM_13)) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~54_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_13),
	.datac(\ALUSrc2_ID~54_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~55_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~55 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N2
cycloneive_lcell_comb \ALUSrc1_ID~38 (
// Equation(s):
// \ALUSrc1_ID~38_combout  = (Instr_IF_25 & (rfifrdat1_13)) # (!Instr_IF_25 & ((rfifrdat1_131)))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_13),
	.datad(rfifrdat1_131),
	.cin(gnd),
	.combout(\ALUSrc1_ID~38_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~38 .lut_mask = 16'hF3C0;
defparam \ALUSrc1_ID~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N16
cycloneive_lcell_comb \ALUSrc1_ID~39 (
// Equation(s):
// \ALUSrc1_ID~39_combout  = (ReadData_MEM_13 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~38_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_13 & (\ALUSrc1_ID~38_combout  & ((\ALUSrc1_ID~1_combout ))))

	.dataa(ReadData_MEM_13),
	.datab(\ALUSrc1_ID~38_combout ),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~39_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~39 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \ALUSrc2_ID~56 (
// Equation(s):
// \ALUSrc2_ID~56_combout  = (Instr_IF[12] & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_12)))) # (!Instr_IF[12] & (((\Equal0~0_combout  & rfifrdat2_12))))

	.dataa(Instr_IF[12]),
	.datab(\ALUSrc2_ID~49_combout ),
	.datac(Equal0),
	.datad(rfifrdat2_12),
	.cin(gnd),
	.combout(\ALUSrc2_ID~56_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~56 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N4
cycloneive_lcell_comb \ALUSrc2_ID~57 (
// Equation(s):
// \ALUSrc2_ID~57_combout  = (\Equal3~0_combout  & (ReadData_MEM_12)) # (!\Equal3~0_combout  & (((!\branch~0_combout  & \ALUSrc2_ID~56_combout ))))

	.dataa(ReadData_MEM_12),
	.datab(branch),
	.datac(\Equal3~0_combout ),
	.datad(\ALUSrc2_ID~56_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~57_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~57 .lut_mask = 16'hA3A0;
defparam \ALUSrc2_ID~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \ALUSrc1_ID~40 (
// Equation(s):
// \ALUSrc1_ID~40_combout  = (Instr_IF_25 & (rfifrdat1_12)) # (!Instr_IF_25 & ((rfifrdat1_121)))

	.dataa(rfifrdat1_12),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_121),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc1_ID~40_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~40 .lut_mask = 16'hB8B8;
defparam \ALUSrc1_ID~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N14
cycloneive_lcell_comb \ALUSrc1_ID~41 (
// Equation(s):
// \ALUSrc1_ID~41_combout  = (ReadData_MEM_12 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~40_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_12 & (\ALUSrc1_ID~40_combout  & ((\ALUSrc1_ID~1_combout ))))

	.dataa(ReadData_MEM_12),
	.datab(\ALUSrc1_ID~40_combout ),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~41_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~41 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N24
cycloneive_lcell_comb \CalcData_MEM[11]~feeder (
// Equation(s):
// \CalcData_MEM[11]~feeder_combout  = Result_EX_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_11),
	.cin(gnd),
	.combout(\CalcData_MEM[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[11]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \ALUSrc2_ID~58 (
// Equation(s):
// \ALUSrc2_ID~58_combout  = (\ALUSrc2_ID~49_combout  & ((Instr_IF[11]) # ((\Equal0~0_combout  & rfifrdat2_11)))) # (!\ALUSrc2_ID~49_combout  & (\Equal0~0_combout  & ((rfifrdat2_11))))

	.dataa(\ALUSrc2_ID~49_combout ),
	.datab(Equal0),
	.datac(Instr_IF[11]),
	.datad(rfifrdat2_11),
	.cin(gnd),
	.combout(\ALUSrc2_ID~58_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~58 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N30
cycloneive_lcell_comb \ALUSrc2_ID~59 (
// Equation(s):
// \ALUSrc2_ID~59_combout  = (\Equal3~0_combout  & (((ReadData_MEM_11)))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~58_combout  & ((!\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(\ALUSrc2_ID~58_combout ),
	.datac(ReadData_MEM_11),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~59_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~59 .lut_mask = 16'hA0E4;
defparam \ALUSrc2_ID~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N18
cycloneive_lcell_comb \ALUSrc1_ID~42 (
// Equation(s):
// \ALUSrc1_ID~42_combout  = (Instr_IF_25 & (rfifrdat1_11)) # (!Instr_IF_25 & ((rfifrdat1_111)))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_11),
	.datad(rfifrdat1_111),
	.cin(gnd),
	.combout(\ALUSrc1_ID~42_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~42 .lut_mask = 16'hF3C0;
defparam \ALUSrc1_ID~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N20
cycloneive_lcell_comb \ALUSrc1_ID~43 (
// Equation(s):
// \ALUSrc1_ID~43_combout  = (\ALUSrc1_ID~42_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_11 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~42_combout  & (ReadData_MEM_11 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~42_combout ),
	.datab(ReadData_MEM_11),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~43_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~43 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N28
cycloneive_lcell_comb \ReadData_MEM[10]~feeder (
// Equation(s):
// \ReadData_MEM[10]~feeder_combout  = ramiframload_10

	.dataa(ramiframload_10),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[10]~feeder .lut_mask = 16'hAAAA;
defparam \ReadData_MEM[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \ALUSrc2_ID~60 (
// Equation(s):
// \ALUSrc2_ID~60_combout  = (Instr_IF_10 & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_10)))) # (!Instr_IF_10 & (\Equal0~0_combout  & ((rfifrdat2_10))))

	.dataa(Instr_IF_10),
	.datab(Equal0),
	.datac(\ALUSrc2_ID~49_combout ),
	.datad(rfifrdat2_10),
	.cin(gnd),
	.combout(\ALUSrc2_ID~60_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~60 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N16
cycloneive_lcell_comb \ALUSrc2_ID~61 (
// Equation(s):
// \ALUSrc2_ID~61_combout  = (\Equal3~0_combout  & (((ReadData_MEM_10)))) # (!\Equal3~0_combout  & (!\branch~0_combout  & ((\ALUSrc2_ID~60_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(branch),
	.datac(ReadData_MEM_10),
	.datad(\ALUSrc2_ID~60_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~61_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~61 .lut_mask = 16'hB1A0;
defparam \ALUSrc2_ID~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N26
cycloneive_lcell_comb \ALUSrc1_ID~44 (
// Equation(s):
// \ALUSrc1_ID~44_combout  = (Instr_IF_25 & ((rfifrdat1_10))) # (!Instr_IF_25 & (rfifrdat1_101))

	.dataa(gnd),
	.datab(rfifrdat1_101),
	.datac(Instr_IF_25),
	.datad(rfifrdat1_10),
	.cin(gnd),
	.combout(\ALUSrc1_ID~44_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~44 .lut_mask = 16'hFC0C;
defparam \ALUSrc1_ID~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N28
cycloneive_lcell_comb \ALUSrc1_ID~45 (
// Equation(s):
// \ALUSrc1_ID~45_combout  = (\Equal20~0_combout  & ((ReadData_MEM_10) # ((\ALUSrc1_ID~44_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~44_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_10),
	.datac(\ALUSrc1_ID~44_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~45_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~45 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \ReadData_MEM[9]~feeder (
// Equation(s):
// \ReadData_MEM[9]~feeder_combout  = ramiframload_9

	.dataa(gnd),
	.datab(ramiframload_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[9]~feeder .lut_mask = 16'hCCCC;
defparam \ReadData_MEM[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \CalcData_MEM[9]~feeder (
// Equation(s):
// \CalcData_MEM[9]~feeder_combout  = Result_EX_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_9),
	.cin(gnd),
	.combout(\CalcData_MEM[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[9]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \ALUSrc2_ID~62 (
// Equation(s):
// \ALUSrc2_ID~62_combout  = (\ALUSrc2_ID~49_combout  & ((Instr_IF_9) # ((rfifrdat2_9 & \Equal0~0_combout )))) # (!\ALUSrc2_ID~49_combout  & (rfifrdat2_9 & (\Equal0~0_combout )))

	.dataa(\ALUSrc2_ID~49_combout ),
	.datab(rfifrdat2_9),
	.datac(Equal0),
	.datad(Instr_IF_9),
	.cin(gnd),
	.combout(\ALUSrc2_ID~62_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~62 .lut_mask = 16'hEAC0;
defparam \ALUSrc2_ID~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \ALUSrc2_ID~63 (
// Equation(s):
// \ALUSrc2_ID~63_combout  = (\Equal3~0_combout  & (((ReadData_MEM_9)))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~62_combout  & (!\branch~0_combout )))

	.dataa(\ALUSrc2_ID~62_combout ),
	.datab(branch),
	.datac(\Equal3~0_combout ),
	.datad(ReadData_MEM_9),
	.cin(gnd),
	.combout(\ALUSrc2_ID~63_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~63 .lut_mask = 16'hF202;
defparam \ALUSrc2_ID~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \ALUSrc1_ID~46 (
// Equation(s):
// \ALUSrc1_ID~46_combout  = (Instr_IF_25 & (rfifrdat1_9)) # (!Instr_IF_25 & ((rfifrdat1_91)))

	.dataa(rfifrdat1_9),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_91),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSrc1_ID~46_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~46 .lut_mask = 16'hB8B8;
defparam \ALUSrc1_ID~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \ALUSrc1_ID~47 (
// Equation(s):
// \ALUSrc1_ID~47_combout  = (\Equal20~0_combout  & ((ReadData_MEM_9) # ((\ALUSrc1_ID~46_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (\ALUSrc1_ID~46_combout  & ((\ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(\ALUSrc1_ID~46_combout ),
	.datac(ReadData_MEM_9),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~47_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~47 .lut_mask = 16'hECA0;
defparam \ALUSrc1_ID~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \ReadData_MEM[8]~feeder (
// Equation(s):
// \ReadData_MEM[8]~feeder_combout  = ramiframload_8

	.dataa(gnd),
	.datab(ramiframload_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[8]~feeder .lut_mask = 16'hCCCC;
defparam \ReadData_MEM[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \ALUSrc2_ID~64 (
// Equation(s):
// \ALUSrc2_ID~64_combout  = (Instr_IF_8 & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_8)))) # (!Instr_IF_8 & (\Equal0~0_combout  & ((rfifrdat2_8))))

	.dataa(Instr_IF_8),
	.datab(Equal0),
	.datac(\ALUSrc2_ID~49_combout ),
	.datad(rfifrdat2_8),
	.cin(gnd),
	.combout(\ALUSrc2_ID~64_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~64 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \ALUSrc2_ID~65 (
// Equation(s):
// \ALUSrc2_ID~65_combout  = (\Equal3~0_combout  & (ReadData_MEM_8)) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~64_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_8),
	.datac(\ALUSrc2_ID~64_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~65_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~65 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \ALUSrc1_ID~48 (
// Equation(s):
// \ALUSrc1_ID~48_combout  = (Instr_IF_25 & (rfifrdat1_8)) # (!Instr_IF_25 & ((rfifrdat1_81)))

	.dataa(rfifrdat1_8),
	.datab(Instr_IF_25),
	.datac(gnd),
	.datad(rfifrdat1_81),
	.cin(gnd),
	.combout(\ALUSrc1_ID~48_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~48 .lut_mask = 16'hBB88;
defparam \ALUSrc1_ID~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \ALUSrc1_ID~49 (
// Equation(s):
// \ALUSrc1_ID~49_combout  = (\Equal20~0_combout  & ((ReadData_MEM_8) # ((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~48_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~48_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_8),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(\ALUSrc1_ID~48_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~49_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~49 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \CalcData_MEM[7]~feeder (
// Equation(s):
// \CalcData_MEM[7]~feeder_combout  = Result_EX_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Result_EX_7),
	.cin(gnd),
	.combout(\CalcData_MEM[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \CalcData_MEM[7]~feeder .lut_mask = 16'hFF00;
defparam \CalcData_MEM[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \ALUSrc2_ID~66 (
// Equation(s):
// \ALUSrc2_ID~66_combout  = (Instr_IF_7 & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_7)))) # (!Instr_IF_7 & (\Equal0~0_combout  & ((rfifrdat2_7))))

	.dataa(Instr_IF_7),
	.datab(Equal0),
	.datac(\ALUSrc2_ID~49_combout ),
	.datad(rfifrdat2_7),
	.cin(gnd),
	.combout(\ALUSrc2_ID~66_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~66 .lut_mask = 16'hECA0;
defparam \ALUSrc2_ID~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \ALUSrc2_ID~67 (
// Equation(s):
// \ALUSrc2_ID~67_combout  = (\Equal3~0_combout  & (ReadData_MEM_7)) # (!\Equal3~0_combout  & (((\ALUSrc2_ID~66_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_7),
	.datac(\ALUSrc2_ID~66_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~67_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~67 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \ALUSrc1_ID~50 (
// Equation(s):
// \ALUSrc1_ID~50_combout  = (Instr_IF_25 & (rfifrdat1_7)) # (!Instr_IF_25 & ((rfifrdat1_71)))

	.dataa(rfifrdat1_7),
	.datab(gnd),
	.datac(Instr_IF_25),
	.datad(rfifrdat1_71),
	.cin(gnd),
	.combout(\ALUSrc1_ID~50_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~50 .lut_mask = 16'hAFA0;
defparam \ALUSrc1_ID~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \ALUSrc1_ID~51 (
// Equation(s):
// \ALUSrc1_ID~51_combout  = (\Equal20~0_combout  & ((ReadData_MEM_7) # ((\ALUSrc1_ID~50_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~50_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_7),
	.datac(\ALUSrc1_ID~50_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~51_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~51 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \ALUSrc2_ID~68 (
// Equation(s):
// \ALUSrc2_ID~68_combout  = (Instr_IF_6 & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_6)))) # (!Instr_IF_6 & (((\Equal0~0_combout  & rfifrdat2_6))))

	.dataa(Instr_IF_6),
	.datab(\ALUSrc2_ID~49_combout ),
	.datac(Equal0),
	.datad(rfifrdat2_6),
	.cin(gnd),
	.combout(\ALUSrc2_ID~68_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~68 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \ALUSrc2_ID~69 (
// Equation(s):
// \ALUSrc2_ID~69_combout  = (\Equal3~0_combout  & (((ReadData_MEM_6)))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~68_combout  & ((!\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(\ALUSrc2_ID~68_combout ),
	.datac(ReadData_MEM_6),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~69_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~69 .lut_mask = 16'hA0E4;
defparam \ALUSrc2_ID~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N24
cycloneive_lcell_comb \ALUSrc1_ID~52 (
// Equation(s):
// \ALUSrc1_ID~52_combout  = (Instr_IF_25 & ((rfifrdat1_6))) # (!Instr_IF_25 & (rfifrdat1_61))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_61),
	.datad(rfifrdat1_6),
	.cin(gnd),
	.combout(\ALUSrc1_ID~52_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~52 .lut_mask = 16'hFC30;
defparam \ALUSrc1_ID~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N20
cycloneive_lcell_comb \ALUSrc1_ID~53 (
// Equation(s):
// \ALUSrc1_ID~53_combout  = (\Equal20~0_combout  & ((ReadData_MEM_6) # ((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~52_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~52_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_6),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(\ALUSrc1_ID~52_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~53_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~53 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \ALUSrc2_ID~70 (
// Equation(s):
// \ALUSrc2_ID~70_combout  = (Instr_IF_5 & ((\ALUSrc2_ID~49_combout ) # ((\Equal0~0_combout  & rfifrdat2_5)))) # (!Instr_IF_5 & (((\Equal0~0_combout  & rfifrdat2_5))))

	.dataa(Instr_IF_5),
	.datab(\ALUSrc2_ID~49_combout ),
	.datac(Equal0),
	.datad(rfifrdat2_5),
	.cin(gnd),
	.combout(\ALUSrc2_ID~70_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~70 .lut_mask = 16'hF888;
defparam \ALUSrc2_ID~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \ALUSrc2_ID~71 (
// Equation(s):
// \ALUSrc2_ID~71_combout  = (\Equal3~0_combout  & (((ReadData_MEM_5)))) # (!\Equal3~0_combout  & (\ALUSrc2_ID~70_combout  & ((!\branch~0_combout ))))

	.dataa(\ALUSrc2_ID~70_combout ),
	.datab(ReadData_MEM_5),
	.datac(branch),
	.datad(\Equal3~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc2_ID~71_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~71 .lut_mask = 16'hCC0A;
defparam \ALUSrc2_ID~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N12
cycloneive_lcell_comb \ALUSrc1_ID~54 (
// Equation(s):
// \ALUSrc1_ID~54_combout  = (Instr_IF_25 & ((rfifrdat1_5))) # (!Instr_IF_25 & (rfifrdat1_51))

	.dataa(rfifrdat1_51),
	.datab(Instr_IF_25),
	.datac(gnd),
	.datad(rfifrdat1_5),
	.cin(gnd),
	.combout(\ALUSrc1_ID~54_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~54 .lut_mask = 16'hEE22;
defparam \ALUSrc1_ID~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N10
cycloneive_lcell_comb \ALUSrc1_ID~55 (
// Equation(s):
// \ALUSrc1_ID~55_combout  = (\Equal20~0_combout  & ((ReadData_MEM_5) # ((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~54_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~54_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_5),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(\ALUSrc1_ID~54_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~55_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~55 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N28
cycloneive_lcell_comb \ReadData_MEM[4]~feeder (
// Equation(s):
// \ReadData_MEM[4]~feeder_combout  = ramiframload_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(\ReadData_MEM[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[4]~feeder .lut_mask = 16'hFF00;
defparam \ReadData_MEM[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N2
cycloneive_lcell_comb \ALUSrc2_ID~72 (
// Equation(s):
// \ALUSrc2_ID~72_combout  = (\Equal3~0_combout  & (((ReadData_MEM_4)))) # (!\Equal3~0_combout  & (!\branch~0_combout  & ((\input_ALUSrc2_ID~3_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(branch),
	.datac(ReadData_MEM_4),
	.datad(input_ALUSrc2_ID),
	.cin(gnd),
	.combout(\ALUSrc2_ID~72_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~72 .lut_mask = 16'hB1A0;
defparam \ALUSrc2_ID~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \ALUSrc1_ID~56 (
// Equation(s):
// \ALUSrc1_ID~56_combout  = (Instr_IF_25 & (rfifrdat1_4)) # (!Instr_IF_25 & ((rfifrdat1_41)))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_4),
	.datac(gnd),
	.datad(rfifrdat1_41),
	.cin(gnd),
	.combout(\ALUSrc1_ID~56_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~56 .lut_mask = 16'hDD88;
defparam \ALUSrc1_ID~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \ALUSrc1_ID~57 (
// Equation(s):
// \ALUSrc1_ID~57_combout  = (\Equal20~0_combout  & ((ReadData_MEM_4) # ((\ALUSrc1_ID~56_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~56_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_4),
	.datac(\ALUSrc1_ID~56_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~57_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~57 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \ALUSrc2_ID~73 (
// Equation(s):
// \ALUSrc2_ID~73_combout  = (\Equal3~0_combout  & (ReadData_MEM_3)) # (!\Equal3~0_combout  & (((\input_ALUSrc2_ID~5_combout  & !\branch~0_combout ))))

	.dataa(ReadData_MEM_3),
	.datab(\Equal3~0_combout ),
	.datac(input_ALUSrc2_ID1),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~73_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~73 .lut_mask = 16'h88B8;
defparam \ALUSrc2_ID~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \ALUSrc1_ID~58 (
// Equation(s):
// \ALUSrc1_ID~58_combout  = (Instr_IF_25 & ((rfifrdat1_3))) # (!Instr_IF_25 & (rfifrdat1_32))

	.dataa(gnd),
	.datab(rfifrdat1_32),
	.datac(Instr_IF_25),
	.datad(rfifrdat1_3),
	.cin(gnd),
	.combout(\ALUSrc1_ID~58_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~58 .lut_mask = 16'hFC0C;
defparam \ALUSrc1_ID~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N0
cycloneive_lcell_comb \ALUSrc1_ID~59 (
// Equation(s):
// \ALUSrc1_ID~59_combout  = (\Equal20~0_combout  & ((ReadData_MEM_3) # ((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~58_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~1_combout  & \ALUSrc1_ID~58_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_3),
	.datac(\ALUSrc1_ID~1_combout ),
	.datad(\ALUSrc1_ID~58_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~59_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~59 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \ALUSrc2_ID~74 (
// Equation(s):
// \ALUSrc2_ID~74_combout  = (\Equal3~0_combout  & (ReadData_MEM_2)) # (!\Equal3~0_combout  & (((\input_ALUSrc2_ID~7_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_2),
	.datac(input_ALUSrc2_ID2),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~74_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~74 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \ALUSrc1_ID~60 (
// Equation(s):
// \ALUSrc1_ID~60_combout  = (Instr_IF_25 & ((rfifrdat1_2))) # (!Instr_IF_25 & (rfifrdat1_210))

	.dataa(Instr_IF_25),
	.datab(rfifrdat1_210),
	.datac(gnd),
	.datad(rfifrdat1_2),
	.cin(gnd),
	.combout(\ALUSrc1_ID~60_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~60 .lut_mask = 16'hEE44;
defparam \ALUSrc1_ID~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \ALUSrc1_ID~61 (
// Equation(s):
// \ALUSrc1_ID~61_combout  = (ReadData_MEM_2 & ((\Equal20~0_combout ) # ((\ALUSrc1_ID~60_combout  & \ALUSrc1_ID~1_combout )))) # (!ReadData_MEM_2 & (((\ALUSrc1_ID~60_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(ReadData_MEM_2),
	.datab(Equal20),
	.datac(\ALUSrc1_ID~60_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~61_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~61 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \ReadData_MEM[1]~feeder (
// Equation(s):
// \ReadData_MEM[1]~feeder_combout  = ramiframload_1

	.dataa(gnd),
	.datab(ramiframload_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ReadData_MEM[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ReadData_MEM[1]~feeder .lut_mask = 16'hCCCC;
defparam \ReadData_MEM[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \ALUSrc2_ID~75 (
// Equation(s):
// \ALUSrc2_ID~75_combout  = (\Equal3~0_combout  & (ReadData_MEM_1)) # (!\Equal3~0_combout  & (((\input_ALUSrc2_ID~9_combout  & !\branch~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(ReadData_MEM_1),
	.datac(input_ALUSrc2_ID3),
	.datad(branch),
	.cin(gnd),
	.combout(\ALUSrc2_ID~75_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~75 .lut_mask = 16'h88D8;
defparam \ALUSrc2_ID~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \ALUSrc1_ID~62 (
// Equation(s):
// \ALUSrc1_ID~62_combout  = (Instr_IF_25 & ((rfifrdat1_1))) # (!Instr_IF_25 & (rfifrdat1_110))

	.dataa(rfifrdat1_110),
	.datab(gnd),
	.datac(Instr_IF_25),
	.datad(rfifrdat1_1),
	.cin(gnd),
	.combout(\ALUSrc1_ID~62_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~62 .lut_mask = 16'hFA0A;
defparam \ALUSrc1_ID~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N6
cycloneive_lcell_comb \ALUSrc1_ID~63 (
// Equation(s):
// \ALUSrc1_ID~63_combout  = (\ALUSrc1_ID~62_combout  & ((\ALUSrc1_ID~1_combout ) # ((ReadData_MEM_1 & \Equal20~0_combout )))) # (!\ALUSrc1_ID~62_combout  & (ReadData_MEM_1 & (\Equal20~0_combout )))

	.dataa(\ALUSrc1_ID~62_combout ),
	.datab(ReadData_MEM_1),
	.datac(Equal20),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~63_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~63 .lut_mask = 16'hEAC0;
defparam \ALUSrc1_ID~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \ALUSrc2_ID~76 (
// Equation(s):
// \ALUSrc2_ID~76_combout  = (\Equal3~0_combout  & (((ReadData_MEM_0)))) # (!\Equal3~0_combout  & (!\branch~0_combout  & ((\input_ALUSrc2_ID~11_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(branch),
	.datac(ReadData_MEM_0),
	.datad(input_ALUSrc2_ID4),
	.cin(gnd),
	.combout(\ALUSrc2_ID~76_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc2_ID~76 .lut_mask = 16'hB1A0;
defparam \ALUSrc2_ID~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \ALUSrc1_ID~64 (
// Equation(s):
// \ALUSrc1_ID~64_combout  = (Instr_IF_25 & (rfifrdat1_0)) # (!Instr_IF_25 & ((rfifrdat1_01)))

	.dataa(gnd),
	.datab(Instr_IF_25),
	.datac(rfifrdat1_0),
	.datad(rfifrdat1_01),
	.cin(gnd),
	.combout(\ALUSrc1_ID~64_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~64 .lut_mask = 16'hF3C0;
defparam \ALUSrc1_ID~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N26
cycloneive_lcell_comb \ALUSrc1_ID~65 (
// Equation(s):
// \ALUSrc1_ID~65_combout  = (\Equal20~0_combout  & ((ReadData_MEM_0) # ((\ALUSrc1_ID~64_combout  & \ALUSrc1_ID~1_combout )))) # (!\Equal20~0_combout  & (((\ALUSrc1_ID~64_combout  & \ALUSrc1_ID~1_combout ))))

	.dataa(Equal20),
	.datab(ReadData_MEM_0),
	.datac(\ALUSrc1_ID~64_combout ),
	.datad(\ALUSrc1_ID~1_combout ),
	.cin(gnd),
	.combout(\ALUSrc1_ID~65_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc1_ID~65 .lut_mask = 16'hF888;
defparam \ALUSrc1_ID~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \Wdata_EX~1 (
// Equation(s):
// \Wdata_EX~1_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_0))) # (!always01 & (RegDat2_ID[0]))))

	.dataa(RegDat2_ID[0]),
	.datab(src2_hazard_t),
	.datac(Result_EX_0),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~1 .lut_mask = 16'h3022;
defparam \Wdata_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \Wdata_EX~0 (
// Equation(s):
// \Wdata_EX~0_combout  = (\always1~0_combout  & (!src2_hazard_t2 & ((!always01) # (!src2_hazard_t1))))

	.dataa(\always1~0_combout ),
	.datab(src2_hazard_t),
	.datac(always0),
	.datad(src2_hazard_t1),
	.cin(gnd),
	.combout(\Wdata_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~0 .lut_mask = 16'h002A;
defparam \Wdata_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \Wdata_EX~2 (
// Equation(s):
// \Wdata_EX~2_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~1_combout ) # ((\input_a~135_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~1_combout ),
	.datab(\Wdata_EX~0_combout ),
	.datac(input_a14),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~2 .lut_mask = 16'hC888;
defparam \Wdata_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \nextPC_IF~0 (
// Equation(s):
// \nextPC_IF~0_combout  = (pc_1 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_1),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~0_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~0 .lut_mask = 16'h00F0;
defparam \nextPC_IF~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N1
dffeas \nextPC_IF[1] (
	.clk(CLK),
	.d(\nextPC_IF~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[1]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[1] .is_wysiwyg = "true";
defparam \nextPC_IF[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \nextPC_ID~0 (
// Equation(s):
// \nextPC_ID~0_combout  = (nextPC_IF[1] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[1]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~0 .lut_mask = 16'h00CC;
defparam \nextPC_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N8
cycloneive_lcell_comb \jump_ID~0 (
// Equation(s):
// \jump_ID~0_combout  = (!Instr_IF_30 & (!Instr_IF_31 & (!\branch~0_combout  & WideOr33)))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_31),
	.datac(branch),
	.datad(WideOr33),
	.cin(gnd),
	.combout(\jump_ID~0_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~0 .lut_mask = 16'h0100;
defparam \jump_ID~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N22
cycloneive_lcell_comb \jump_ID~1 (
// Equation(s):
// \jump_ID~1_combout  = (!Instr_IF_30 & (!Instr_IF_26 & (!Instr_IF_29 & Instr_IF_28)))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_26),
	.datac(Instr_IF_29),
	.datad(Instr_IF_28),
	.cin(gnd),
	.combout(\jump_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~1 .lut_mask = 16'h0100;
defparam \jump_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N28
cycloneive_lcell_comb \jump_ID~2 (
// Equation(s):
// \jump_ID~2_combout  = (!\branch~0_combout  & ((\jump_ID~1_combout ) # ((Decoder0 & !Selector11))))

	.dataa(\jump_ID~1_combout ),
	.datab(Decoder0),
	.datac(Selector111),
	.datad(branch),
	.cin(gnd),
	.combout(\jump_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~2 .lut_mask = 16'h00AE;
defparam \jump_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \jump_ID~3 (
// Equation(s):
// \jump_ID~3_combout  = (Instr_IF_28 & (!Instr_IF_31 & (!Instr_IF_27 & !Instr_IF_29)))

	.dataa(Instr_IF_28),
	.datab(Instr_IF_31),
	.datac(Instr_IF_27),
	.datad(Instr_IF_29),
	.cin(gnd),
	.combout(\jump_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~3 .lut_mask = 16'h0002;
defparam \jump_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \jump_ID~4 (
// Equation(s):
// \jump_ID~4_combout  = (!Instr_IF_30 & (Instr_IF_26 & (\jump_ID~3_combout  & !\branch~0_combout )))

	.dataa(Instr_IF_30),
	.datab(Instr_IF_26),
	.datac(\jump_ID~3_combout ),
	.datad(branch),
	.cin(gnd),
	.combout(\jump_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \jump_ID~4 .lut_mask = 16'h0040;
defparam \jump_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \nextPC_IF~1 (
// Equation(s):
// \nextPC_IF~1_combout  = (pc_0 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_0),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~1_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~1 .lut_mask = 16'h00F0;
defparam \nextPC_IF~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N3
dffeas \nextPC_IF[0] (
	.clk(CLK),
	.d(\nextPC_IF~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[0]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[0] .is_wysiwyg = "true";
defparam \nextPC_IF[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \nextPC_ID~1 (
// Equation(s):
// \nextPC_ID~1_combout  = (nextPC_IF[0] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[0]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~1 .lut_mask = 16'h00CC;
defparam \nextPC_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \nextPC_IF~2 (
// Equation(s):
// \nextPC_IF~2_combout  = (!\branch~0_combout  & \pc_next_plus4[3]~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_3),
	.cin(gnd),
	.combout(\nextPC_IF~2_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~2 .lut_mask = 16'h0F00;
defparam \nextPC_IF~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N3
dffeas \nextPC_IF[3] (
	.clk(CLK),
	.d(\nextPC_IF~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[3]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[3] .is_wysiwyg = "true";
defparam \nextPC_IF[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \nextPC_ID~2 (
// Equation(s):
// \nextPC_ID~2_combout  = (!\branch~0_combout  & nextPC_IF[3])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[3]),
	.cin(gnd),
	.combout(\nextPC_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~2 .lut_mask = 16'h0F00;
defparam \nextPC_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \Instr_ID~10 (
// Equation(s):
// \Instr_ID~10_combout  = (Instr_IF_1 & !\branch~0_combout )

	.dataa(Instr_IF_1),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~10 .lut_mask = 16'h0A0A;
defparam \Instr_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \nextPC_IF~3 (
// Equation(s):
// \nextPC_IF~3_combout  = (!\branch~0_combout  & \pc_next_plus4[2]~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_2),
	.cin(gnd),
	.combout(\nextPC_IF~3_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~3 .lut_mask = 16'h0F00;
defparam \nextPC_IF~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N21
dffeas \nextPC_IF[2] (
	.clk(CLK),
	.d(\nextPC_IF~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[2]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[2] .is_wysiwyg = "true";
defparam \nextPC_IF[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \nextPC_ID~3 (
// Equation(s):
// \nextPC_ID~3_combout  = (!\branch~0_combout  & nextPC_IF[2])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[2]),
	.cin(gnd),
	.combout(\nextPC_ID~3_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~3 .lut_mask = 16'h0F00;
defparam \nextPC_ID~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \Instr_ID~11 (
// Equation(s):
// \Instr_ID~11_combout  = (Instr_IF_0 & !\branch~0_combout )

	.dataa(Instr_IF_0),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~11 .lut_mask = 16'h0A0A;
defparam \Instr_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \nextPC_IF~4 (
// Equation(s):
// \nextPC_IF~4_combout  = (\pc_next_plus4[5]~6_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_5),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~4_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~4 .lut_mask = 16'h00CC;
defparam \nextPC_IF~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N25
dffeas \nextPC_IF[5] (
	.clk(CLK),
	.d(\nextPC_IF~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[5]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[5] .is_wysiwyg = "true";
defparam \nextPC_IF[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \nextPC_ID~4 (
// Equation(s):
// \nextPC_ID~4_combout  = (nextPC_IF[5] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[5]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~4_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~4 .lut_mask = 16'h00CC;
defparam \nextPC_ID~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Instr_ID~12 (
// Equation(s):
// \Instr_ID~12_combout  = (Instr_IF_3 & !\branch~0_combout )

	.dataa(Instr_IF_3),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~12 .lut_mask = 16'h00AA;
defparam \Instr_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \nextPC_IF~5 (
// Equation(s):
// \nextPC_IF~5_combout  = (\pc_next_plus4[4]~4_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_next_plus4_4),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~5_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~5 .lut_mask = 16'h00F0;
defparam \nextPC_IF~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \nextPC_IF[4] (
	.clk(CLK),
	.d(\nextPC_IF~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[4]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[4] .is_wysiwyg = "true";
defparam \nextPC_IF[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \nextPC_ID~5 (
// Equation(s):
// \nextPC_ID~5_combout  = (nextPC_IF[4] & !\branch~0_combout )

	.dataa(nextPC_IF[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~5 .lut_mask = 16'h00AA;
defparam \nextPC_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \Instr_ID~13 (
// Equation(s):
// \Instr_ID~13_combout  = (Instr_IF_2 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_2),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~13 .lut_mask = 16'h00CC;
defparam \Instr_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \nextPC_IF~6 (
// Equation(s):
// \nextPC_IF~6_combout  = (\pc_next_plus4[7]~10_combout  & !\branch~0_combout )

	.dataa(pc_next_plus4_7),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~6_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~6 .lut_mask = 16'h00AA;
defparam \nextPC_IF~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N15
dffeas \nextPC_IF[7] (
	.clk(CLK),
	.d(\nextPC_IF~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[7]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[7] .is_wysiwyg = "true";
defparam \nextPC_IF[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \nextPC_ID~6 (
// Equation(s):
// \nextPC_ID~6_combout  = (nextPC_IF[7] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[7]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~6 .lut_mask = 16'h00CC;
defparam \nextPC_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \Instr_ID~14 (
// Equation(s):
// \Instr_ID~14_combout  = (Instr_IF_5 & !\branch~0_combout )

	.dataa(Instr_IF_5),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~14 .lut_mask = 16'h0A0A;
defparam \Instr_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \nextPC_IF~7 (
// Equation(s):
// \nextPC_IF~7_combout  = (\pc_next_plus4[6]~8_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_next_plus4_6),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~7_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~7 .lut_mask = 16'h00F0;
defparam \nextPC_IF~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N25
dffeas \nextPC_IF[6] (
	.clk(CLK),
	.d(\nextPC_IF~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[6]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[6] .is_wysiwyg = "true";
defparam \nextPC_IF[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \nextPC_ID~7 (
// Equation(s):
// \nextPC_ID~7_combout  = (nextPC_IF[6] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[6]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~7 .lut_mask = 16'h00CC;
defparam \nextPC_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \Instr_ID~15 (
// Equation(s):
// \Instr_ID~15_combout  = (!\branch~0_combout  & Instr_IF_4)

	.dataa(gnd),
	.datab(branch),
	.datac(Instr_IF_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~15 .lut_mask = 16'h3030;
defparam \Instr_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N14
cycloneive_lcell_comb \nextPC_IF~8 (
// Equation(s):
// \nextPC_IF~8_combout  = (!\branch~0_combout  & \pc_next_plus4[9]~14_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_9),
	.cin(gnd),
	.combout(\nextPC_IF~8_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~8 .lut_mask = 16'h0F00;
defparam \nextPC_IF~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N15
dffeas \nextPC_IF[9] (
	.clk(CLK),
	.d(\nextPC_IF~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[9]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[9] .is_wysiwyg = "true";
defparam \nextPC_IF[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N14
cycloneive_lcell_comb \nextPC_ID~8 (
// Equation(s):
// \nextPC_ID~8_combout  = (!\branch~0_combout  & nextPC_IF[9])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[9]),
	.cin(gnd),
	.combout(\nextPC_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~8 .lut_mask = 16'h0F00;
defparam \nextPC_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \Instr_ID~16 (
// Equation(s):
// \Instr_ID~16_combout  = (!\branch~0_combout  & Instr_IF_7)

	.dataa(gnd),
	.datab(branch),
	.datac(Instr_IF_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~16 .lut_mask = 16'h3030;
defparam \Instr_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \nextPC_IF~9 (
// Equation(s):
// \nextPC_IF~9_combout  = (\pc_next_plus4[8]~12_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_8),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~9_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~9 .lut_mask = 16'h00CC;
defparam \nextPC_IF~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N27
dffeas \nextPC_IF[8] (
	.clk(CLK),
	.d(\nextPC_IF~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[8]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[8] .is_wysiwyg = "true";
defparam \nextPC_IF[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \nextPC_ID~9 (
// Equation(s):
// \nextPC_ID~9_combout  = (nextPC_IF[8] & !\branch~0_combout )

	.dataa(nextPC_IF[8]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~9 .lut_mask = 16'h00AA;
defparam \nextPC_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \Instr_ID~17 (
// Equation(s):
// \Instr_ID~17_combout  = (Instr_IF_6 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_6),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~17_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~17 .lut_mask = 16'h00CC;
defparam \Instr_ID~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \nextPC_IF~10 (
// Equation(s):
// \nextPC_IF~10_combout  = (\pc_next_plus4[11]~18_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_11),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~10_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~10 .lut_mask = 16'h00CC;
defparam \nextPC_IF~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N23
dffeas \nextPC_IF[11] (
	.clk(CLK),
	.d(\nextPC_IF~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[11]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[11] .is_wysiwyg = "true";
defparam \nextPC_IF[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \nextPC_ID~10 (
// Equation(s):
// \nextPC_ID~10_combout  = (nextPC_IF[11] & !\branch~0_combout )

	.dataa(nextPC_IF[11]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~10 .lut_mask = 16'h00AA;
defparam \nextPC_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \Instr_ID~18 (
// Equation(s):
// \Instr_ID~18_combout  = (Instr_IF_9 & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF_9),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~18_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~18 .lut_mask = 16'h00CC;
defparam \Instr_ID~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \nextPC_IF~11 (
// Equation(s):
// \nextPC_IF~11_combout  = (\pc_next_plus4[10]~16_combout  & !\branch~0_combout )

	.dataa(pc_next_plus4_10),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~11_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~11 .lut_mask = 16'h00AA;
defparam \nextPC_IF~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N5
dffeas \nextPC_IF[10] (
	.clk(CLK),
	.d(\nextPC_IF~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[10]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[10] .is_wysiwyg = "true";
defparam \nextPC_IF[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \nextPC_ID~11 (
// Equation(s):
// \nextPC_ID~11_combout  = (nextPC_IF[10] & !\branch~0_combout )

	.dataa(nextPC_IF[10]),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~11 .lut_mask = 16'h0A0A;
defparam \nextPC_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N0
cycloneive_lcell_comb \Instr_ID~19 (
// Equation(s):
// \Instr_ID~19_combout  = (Instr_IF_8 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Instr_IF_8),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~19_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~19 .lut_mask = 16'h00F0;
defparam \Instr_ID~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \nextPC_IF~12 (
// Equation(s):
// \nextPC_IF~12_combout  = (\pc_next_plus4[13]~22_combout  & !\branch~0_combout )

	.dataa(pc_next_plus4_13),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~12_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~12 .lut_mask = 16'h0A0A;
defparam \nextPC_IF~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N13
dffeas \nextPC_IF[13] (
	.clk(CLK),
	.d(\nextPC_IF~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[13]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[13] .is_wysiwyg = "true";
defparam \nextPC_IF[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \nextPC_ID~12 (
// Equation(s):
// \nextPC_ID~12_combout  = (!\branch~0_combout  & nextPC_IF[13])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[13]),
	.cin(gnd),
	.combout(\nextPC_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~12 .lut_mask = 16'h0F00;
defparam \nextPC_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \Instr_ID~20 (
// Equation(s):
// \Instr_ID~20_combout  = (Instr_IF[11] & !\branch~0_combout )

	.dataa(Instr_IF[11]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~20_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~20 .lut_mask = 16'h00AA;
defparam \Instr_ID~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \nextPC_IF~13 (
// Equation(s):
// \nextPC_IF~13_combout  = (\pc_next_plus4[12]~20_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_12),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~13_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~13 .lut_mask = 16'h00CC;
defparam \nextPC_IF~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N7
dffeas \nextPC_IF[12] (
	.clk(CLK),
	.d(\nextPC_IF~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[12]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[12] .is_wysiwyg = "true";
defparam \nextPC_IF[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \nextPC_ID~13 (
// Equation(s):
// \nextPC_ID~13_combout  = (nextPC_IF[12] & !\branch~0_combout )

	.dataa(nextPC_IF[12]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~13_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~13 .lut_mask = 16'h00AA;
defparam \nextPC_ID~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \Instr_ID~21 (
// Equation(s):
// \Instr_ID~21_combout  = (Instr_IF_10 & !\branch~0_combout )

	.dataa(Instr_IF_10),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~21_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~21 .lut_mask = 16'h0A0A;
defparam \Instr_ID~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \nextPC_IF~14 (
// Equation(s):
// \nextPC_IF~14_combout  = (!\branch~0_combout  & \pc_next_plus4[15]~26_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_15),
	.cin(gnd),
	.combout(\nextPC_IF~14_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~14 .lut_mask = 16'h0F00;
defparam \nextPC_IF~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N23
dffeas \nextPC_IF[15] (
	.clk(CLK),
	.d(\nextPC_IF~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[15]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[15] .is_wysiwyg = "true";
defparam \nextPC_IF[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \nextPC_ID~14 (
// Equation(s):
// \nextPC_ID~14_combout  = (nextPC_IF[15] & !\branch~0_combout )

	.dataa(nextPC_IF[15]),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~14 .lut_mask = 16'h0A0A;
defparam \nextPC_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \Instr_ID~22 (
// Equation(s):
// \Instr_ID~22_combout  = (Instr_IF[13] & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF[13]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~22_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~22 .lut_mask = 16'h00CC;
defparam \Instr_ID~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \nextPC_IF~15 (
// Equation(s):
// \nextPC_IF~15_combout  = (\pc_next_plus4[14]~24_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_14),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~15_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~15 .lut_mask = 16'h00CC;
defparam \nextPC_IF~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N15
dffeas \nextPC_IF[14] (
	.clk(CLK),
	.d(\nextPC_IF~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[14]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[14] .is_wysiwyg = "true";
defparam \nextPC_IF[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \nextPC_ID~15 (
// Equation(s):
// \nextPC_ID~15_combout  = (nextPC_IF[14] & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(nextPC_IF[14]),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~15 .lut_mask = 16'h00F0;
defparam \nextPC_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N30
cycloneive_lcell_comb \Instr_ID~23 (
// Equation(s):
// \Instr_ID~23_combout  = (Instr_IF[12] & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF[12]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_ID~23_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~23 .lut_mask = 16'h00CC;
defparam \Instr_ID~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \nextPC_IF~16 (
// Equation(s):
// \nextPC_IF~16_combout  = (\pc_next_plus4[17]~30_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_17),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~16_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~16 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N27
dffeas \nextPC_IF[17] (
	.clk(CLK),
	.d(\nextPC_IF~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[17]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[17] .is_wysiwyg = "true";
defparam \nextPC_IF[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \nextPC_ID~16 (
// Equation(s):
// \nextPC_ID~16_combout  = (nextPC_IF[17] & !\branch~0_combout )

	.dataa(nextPC_IF[17]),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~16 .lut_mask = 16'h0A0A;
defparam \nextPC_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \Instr_ID~24 (
// Equation(s):
// \Instr_ID~24_combout  = (Instr_IF[15] & !\branch~0_combout )

	.dataa(gnd),
	.datab(Instr_IF[15]),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~24_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~24 .lut_mask = 16'h0C0C;
defparam \Instr_ID~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \nextPC_IF~17 (
// Equation(s):
// \nextPC_IF~17_combout  = (\pc_next_plus4[16]~28_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_16),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~17_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~17 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N29
dffeas \nextPC_IF[16] (
	.clk(CLK),
	.d(\nextPC_IF~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[16]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[16] .is_wysiwyg = "true";
defparam \nextPC_IF[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \nextPC_ID~17 (
// Equation(s):
// \nextPC_ID~17_combout  = (!\branch~0_combout  & nextPC_IF[16])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[16]),
	.cin(gnd),
	.combout(\nextPC_ID~17_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~17 .lut_mask = 16'h0F00;
defparam \nextPC_ID~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \Instr_ID~25 (
// Equation(s):
// \Instr_ID~25_combout  = (Instr_IF[14] & !\branch~0_combout )

	.dataa(Instr_IF[14]),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\Instr_ID~25_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_ID~25 .lut_mask = 16'h0A0A;
defparam \Instr_ID~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N18
cycloneive_lcell_comb \nextPC_IF~18 (
// Equation(s):
// \nextPC_IF~18_combout  = (!\branch~0_combout  & \pc_next_plus4[19]~34_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_19),
	.cin(gnd),
	.combout(\nextPC_IF~18_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~18 .lut_mask = 16'h0F00;
defparam \nextPC_IF~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N19
dffeas \nextPC_IF[19] (
	.clk(CLK),
	.d(\nextPC_IF~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[19]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[19] .is_wysiwyg = "true";
defparam \nextPC_IF[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N6
cycloneive_lcell_comb \nextPC_ID~18 (
// Equation(s):
// \nextPC_ID~18_combout  = (!\branch~0_combout  & nextPC_IF[19])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[19]),
	.cin(gnd),
	.combout(\nextPC_ID~18_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~18 .lut_mask = 16'h0F00;
defparam \nextPC_ID~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \nextPC_IF~19 (
// Equation(s):
// \nextPC_IF~19_combout  = (!\branch~0_combout  & \pc_next_plus4[18]~32_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_18),
	.cin(gnd),
	.combout(\nextPC_IF~19_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~19 .lut_mask = 16'h0F00;
defparam \nextPC_IF~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N3
dffeas \nextPC_IF[18] (
	.clk(CLK),
	.d(\nextPC_IF~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[18]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[18] .is_wysiwyg = "true";
defparam \nextPC_IF[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \nextPC_ID~19 (
// Equation(s):
// \nextPC_ID~19_combout  = (!\branch~0_combout  & nextPC_IF[18])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[18]),
	.cin(gnd),
	.combout(\nextPC_ID~19_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~19 .lut_mask = 16'h0F00;
defparam \nextPC_ID~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N2
cycloneive_lcell_comb \nextPC_IF~20 (
// Equation(s):
// \nextPC_IF~20_combout  = (\pc_next_plus4[21]~38_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_21),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~20_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~20 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N3
dffeas \nextPC_IF[21] (
	.clk(CLK),
	.d(\nextPC_IF~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[21]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[21] .is_wysiwyg = "true";
defparam \nextPC_IF[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N6
cycloneive_lcell_comb \nextPC_ID~20 (
// Equation(s):
// \nextPC_ID~20_combout  = (!\branch~0_combout  & nextPC_IF[21])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[21]),
	.cin(gnd),
	.combout(\nextPC_ID~20_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~20 .lut_mask = 16'h0F00;
defparam \nextPC_ID~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N4
cycloneive_lcell_comb \nextPC_IF~21 (
// Equation(s):
// \nextPC_IF~21_combout  = (!\branch~0_combout  & \pc_next_plus4[20]~36_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_20),
	.cin(gnd),
	.combout(\nextPC_IF~21_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~21 .lut_mask = 16'h0F00;
defparam \nextPC_IF~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N5
dffeas \nextPC_IF[20] (
	.clk(CLK),
	.d(\nextPC_IF~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[20]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[20] .is_wysiwyg = "true";
defparam \nextPC_IF[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N28
cycloneive_lcell_comb \nextPC_ID~21 (
// Equation(s):
// \nextPC_ID~21_combout  = (nextPC_IF[20] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[20]),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~21_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~21 .lut_mask = 16'h0C0C;
defparam \nextPC_ID~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N26
cycloneive_lcell_comb \nextPC_IF~22 (
// Equation(s):
// \nextPC_IF~22_combout  = (\pc_next_plus4[23]~42_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_23),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~22_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~22 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N27
dffeas \nextPC_IF[23] (
	.clk(CLK),
	.d(\nextPC_IF~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[23]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[23] .is_wysiwyg = "true";
defparam \nextPC_IF[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N30
cycloneive_lcell_comb \nextPC_ID~22 (
// Equation(s):
// \nextPC_ID~22_combout  = (nextPC_IF[23] & !\branch~0_combout )

	.dataa(nextPC_IF[23]),
	.datab(gnd),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~22_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~22 .lut_mask = 16'h0A0A;
defparam \nextPC_ID~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N0
cycloneive_lcell_comb \nextPC_IF~23 (
// Equation(s):
// \nextPC_IF~23_combout  = (\pc_next_plus4[22]~40_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_22),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~23_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~23 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N1
dffeas \nextPC_IF[22] (
	.clk(CLK),
	.d(\nextPC_IF~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[22]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[22] .is_wysiwyg = "true";
defparam \nextPC_IF[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N16
cycloneive_lcell_comb \nextPC_ID~23 (
// Equation(s):
// \nextPC_ID~23_combout  = (!\branch~0_combout  & nextPC_IF[22])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[22]),
	.cin(gnd),
	.combout(\nextPC_ID~23_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~23 .lut_mask = 16'h0F00;
defparam \nextPC_ID~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \nextPC_IF~24 (
// Equation(s):
// \nextPC_IF~24_combout  = (\pc_next_plus4[25]~46_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_25),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~24_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~24 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N13
dffeas \nextPC_IF[25] (
	.clk(CLK),
	.d(\nextPC_IF~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[25]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[25] .is_wysiwyg = "true";
defparam \nextPC_IF[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N4
cycloneive_lcell_comb \nextPC_ID~24 (
// Equation(s):
// \nextPC_ID~24_combout  = (!\branch~0_combout  & nextPC_IF[25])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[25]),
	.cin(gnd),
	.combout(\nextPC_ID~24_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~24 .lut_mask = 16'h0F00;
defparam \nextPC_ID~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \nextPC_IF~25 (
// Equation(s):
// \nextPC_IF~25_combout  = (\pc_next_plus4[24]~44_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_24),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~25_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~25 .lut_mask = 16'h00CC;
defparam \nextPC_IF~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N21
dffeas \nextPC_IF[24] (
	.clk(CLK),
	.d(\nextPC_IF~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[24]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[24] .is_wysiwyg = "true";
defparam \nextPC_IF[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \nextPC_ID~25 (
// Equation(s):
// \nextPC_ID~25_combout  = (nextPC_IF[24] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[24]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~25_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~25 .lut_mask = 16'h00CC;
defparam \nextPC_ID~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \nextPC_IF~26 (
// Equation(s):
// \nextPC_IF~26_combout  = (\pc_next_plus4[27]~50_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_next_plus4_27),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~26_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~26 .lut_mask = 16'h00F0;
defparam \nextPC_IF~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N19
dffeas \nextPC_IF[27] (
	.clk(CLK),
	.d(\nextPC_IF~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[27]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[27] .is_wysiwyg = "true";
defparam \nextPC_IF[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \nextPC_ID~26 (
// Equation(s):
// \nextPC_ID~26_combout  = (nextPC_IF[27] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[27]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~26_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~26 .lut_mask = 16'h00CC;
defparam \nextPC_ID~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \nextPC_IF~27 (
// Equation(s):
// \nextPC_IF~27_combout  = (\pc_next_plus4[26]~48_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_26),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_IF~27_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~27 .lut_mask = 16'h0C0C;
defparam \nextPC_IF~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N5
dffeas \nextPC_IF[26] (
	.clk(CLK),
	.d(\nextPC_IF~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[26]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[26] .is_wysiwyg = "true";
defparam \nextPC_IF[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \nextPC_ID~27 (
// Equation(s):
// \nextPC_ID~27_combout  = (nextPC_IF[26] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[26]),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextPC_ID~27_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~27 .lut_mask = 16'h0C0C;
defparam \nextPC_ID~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \nextPC_IF~28 (
// Equation(s):
// \nextPC_IF~28_combout  = (\pc_next_plus4[29]~54_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_next_plus4_29),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~28_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~28 .lut_mask = 16'h00F0;
defparam \nextPC_IF~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N17
dffeas \nextPC_IF[29] (
	.clk(CLK),
	.d(\nextPC_IF~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[29]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[29] .is_wysiwyg = "true";
defparam \nextPC_IF[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \nextPC_ID~28 (
// Equation(s):
// \nextPC_ID~28_combout  = (nextPC_IF[29] & !\branch~0_combout )

	.dataa(gnd),
	.datab(nextPC_IF[29]),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~28_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~28 .lut_mask = 16'h00CC;
defparam \nextPC_ID~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \nextPC_IF~29 (
// Equation(s):
// \nextPC_IF~29_combout  = (\pc_next_plus4[28]~52_combout  & !\branch~0_combout )

	.dataa(gnd),
	.datab(pc_next_plus4_28),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~29_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~29 .lut_mask = 16'h00CC;
defparam \nextPC_IF~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N23
dffeas \nextPC_IF[28] (
	.clk(CLK),
	.d(\nextPC_IF~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[28]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[28] .is_wysiwyg = "true";
defparam \nextPC_IF[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \nextPC_ID~29 (
// Equation(s):
// \nextPC_ID~29_combout  = (nextPC_IF[28] & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(nextPC_IF[28]),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~29_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~29 .lut_mask = 16'h00F0;
defparam \nextPC_ID~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N22
cycloneive_lcell_comb \nextPC_IF~30 (
// Equation(s):
// \nextPC_IF~30_combout  = (!\branch~0_combout  & \pc_next_plus4[31]~58_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(pc_next_plus4_31),
	.cin(gnd),
	.combout(\nextPC_IF~30_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~30 .lut_mask = 16'h0F00;
defparam \nextPC_IF~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N23
dffeas \nextPC_IF[31] (
	.clk(CLK),
	.d(\nextPC_IF~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[31]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[31] .is_wysiwyg = "true";
defparam \nextPC_IF[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \nextPC_ID~30 (
// Equation(s):
// \nextPC_ID~30_combout  = (!\branch~0_combout  & nextPC_IF[31])

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(nextPC_IF[31]),
	.cin(gnd),
	.combout(\nextPC_ID~30_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~30 .lut_mask = 16'h0F00;
defparam \nextPC_ID~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \nextPC_IF~31 (
// Equation(s):
// \nextPC_IF~31_combout  = (\pc_next_plus4[30]~56_combout  & !\branch~0_combout )

	.dataa(pc_next_plus4_30),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_IF~31_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_IF~31 .lut_mask = 16'h00AA;
defparam \nextPC_IF~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N13
dffeas \nextPC_IF[30] (
	.clk(CLK),
	.d(\nextPC_IF~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(nextPC_IF[30]),
	.prn(vcc));
// synopsys translate_off
defparam \nextPC_IF[30] .is_wysiwyg = "true";
defparam \nextPC_IF[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \nextPC_ID~31 (
// Equation(s):
// \nextPC_ID~31_combout  = (nextPC_IF[30] & !\branch~0_combout )

	.dataa(nextPC_IF[30]),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\nextPC_ID~31_combout ),
	.cout());
// synopsys translate_off
defparam \nextPC_ID~31 .lut_mask = 16'h00AA;
defparam \nextPC_ID~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \RegDat2_ID~1 (
// Equation(s):
// \RegDat2_ID~1_combout  = (rfifrdat2_1 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_1),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDat2_ID~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~1 .lut_mask = 16'h0C0C;
defparam \RegDat2_ID~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N17
dffeas \RegDat2_ID[1] (
	.clk(CLK),
	.d(\RegDat2_ID~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[1]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[1] .is_wysiwyg = "true";
defparam \RegDat2_ID[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Wdata_EX~3 (
// Equation(s):
// \Wdata_EX~3_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_1))) # (!always01 & (RegDat2_ID[1]))))

	.dataa(src2_hazard_t),
	.datab(RegDat2_ID[1]),
	.datac(Result_EX_1),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~3 .lut_mask = 16'h5044;
defparam \Wdata_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Wdata_EX~4 (
// Equation(s):
// \Wdata_EX~4_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~3_combout ) # ((\input_a~132_combout  & \Equal27~0_combout ))))

	.dataa(input_a13),
	.datab(\Wdata_EX~3_combout ),
	.datac(\Wdata_EX~0_combout ),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~4 .lut_mask = 16'hE0C0;
defparam \Wdata_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \RegDat2_ID~2 (
// Equation(s):
// \RegDat2_ID~2_combout  = (!\branch~0_combout  & rfifrdat2_2)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_2),
	.cin(gnd),
	.combout(\RegDat2_ID~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~2 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N25
dffeas \RegDat2_ID[2] (
	.clk(CLK),
	.d(\RegDat2_ID~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[2]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[2] .is_wysiwyg = "true";
defparam \RegDat2_ID[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \Wdata_EX~5 (
// Equation(s):
// \Wdata_EX~5_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_2)) # (!always01 & ((RegDat2_ID[2])))))

	.dataa(Result_EX_2),
	.datab(RegDat2_ID[2]),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~5 .lut_mask = 16'h0A0C;
defparam \Wdata_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \Wdata_EX~6 (
// Equation(s):
// \Wdata_EX~6_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~5_combout ) # ((\input_a~129_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(\Wdata_EX~5_combout ),
	.datac(input_a12),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~6 .lut_mask = 16'hA888;
defparam \Wdata_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \Wdata_EX~7 (
// Equation(s):
// \Wdata_EX~7_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_3))) # (!always01 & (RegDat2_ID[3]))))

	.dataa(RegDat2_ID[3]),
	.datab(Result_EX_3),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~7 .lut_mask = 16'h0C0A;
defparam \Wdata_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \Wdata_EX~8 (
// Equation(s):
// \Wdata_EX~8_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~7_combout ) # ((\input_a~126_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~7_combout ),
	.datab(input_a11),
	.datac(Equal27),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~8 .lut_mask = 16'hEA00;
defparam \Wdata_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N0
cycloneive_lcell_comb \Wdata_EX~9 (
// Equation(s):
// \Wdata_EX~9_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_4))) # (!always01 & (RegDat2_ID[4]))))

	.dataa(RegDat2_ID[4]),
	.datab(always0),
	.datac(Result_EX_4),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~9 .lut_mask = 16'h00E2;
defparam \Wdata_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N8
cycloneive_lcell_comb \Wdata_EX~10 (
// Equation(s):
// \Wdata_EX~10_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~9_combout ) # ((\Equal27~0_combout  & \input_a~123_combout ))))

	.dataa(Equal27),
	.datab(input_a10),
	.datac(\Wdata_EX~0_combout ),
	.datad(\Wdata_EX~9_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~10 .lut_mask = 16'hF080;
defparam \Wdata_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \RegDat2_ID~5 (
// Equation(s):
// \RegDat2_ID~5_combout  = (rfifrdat2_5 & !\branch~0_combout )

	.dataa(rfifrdat2_5),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~5_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~5 .lut_mask = 16'h00AA;
defparam \RegDat2_ID~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N29
dffeas \RegDat2_ID[5] (
	.clk(CLK),
	.d(\RegDat2_ID~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[5]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[5] .is_wysiwyg = "true";
defparam \RegDat2_ID[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Wdata_EX~11 (
// Equation(s):
// \Wdata_EX~11_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_5))) # (!always01 & (RegDat2_ID[5]))))

	.dataa(src2_hazard_t),
	.datab(RegDat2_ID[5]),
	.datac(Result_EX_5),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~11 .lut_mask = 16'h5044;
defparam \Wdata_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \Wdata_EX~12 (
// Equation(s):
// \Wdata_EX~12_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~11_combout ) # ((\input_a~120_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~11_combout ),
	.datab(input_a9),
	.datac(Equal27),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~12 .lut_mask = 16'hEA00;
defparam \Wdata_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \RegDat2_ID~6 (
// Equation(s):
// \RegDat2_ID~6_combout  = (rfifrdat2_6 & !\branch~0_combout )

	.dataa(rfifrdat2_6),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~6_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~6 .lut_mask = 16'h00AA;
defparam \RegDat2_ID~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N1
dffeas \RegDat2_ID[6] (
	.clk(CLK),
	.d(\RegDat2_ID~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[6]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[6] .is_wysiwyg = "true";
defparam \RegDat2_ID[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \Wdata_EX~13 (
// Equation(s):
// \Wdata_EX~13_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_6))) # (!always01 & (RegDat2_ID[6]))))

	.dataa(always0),
	.datab(RegDat2_ID[6]),
	.datac(Result_EX_6),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~13 .lut_mask = 16'h00E4;
defparam \Wdata_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \Wdata_EX~14 (
// Equation(s):
// \Wdata_EX~14_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~13_combout ) # ((\Equal27~0_combout  & \input_a~117_combout ))))

	.dataa(Equal27),
	.datab(\Wdata_EX~13_combout ),
	.datac(input_a8),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~14 .lut_mask = 16'hEC00;
defparam \Wdata_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \RegDat2_ID~7 (
// Equation(s):
// \RegDat2_ID~7_combout  = (rfifrdat2_7 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_7),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~7_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~7 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N15
dffeas \RegDat2_ID[7] (
	.clk(CLK),
	.d(\RegDat2_ID~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[7]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[7] .is_wysiwyg = "true";
defparam \RegDat2_ID[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \Wdata_EX~15 (
// Equation(s):
// \Wdata_EX~15_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_7)) # (!always01 & ((RegDat2_ID[7])))))

	.dataa(Result_EX_7),
	.datab(always0),
	.datac(src2_hazard_t),
	.datad(RegDat2_ID[7]),
	.cin(gnd),
	.combout(\Wdata_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~15 .lut_mask = 16'h0B08;
defparam \Wdata_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \Wdata_EX~16 (
// Equation(s):
// \Wdata_EX~16_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~15_combout ) # ((\Equal27~0_combout  & \input_a~114_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(\Wdata_EX~15_combout ),
	.datac(Equal27),
	.datad(input_a7),
	.cin(gnd),
	.combout(\Wdata_EX~16_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~16 .lut_mask = 16'hA888;
defparam \Wdata_EX~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \RegDat2_ID~8 (
// Equation(s):
// \RegDat2_ID~8_combout  = (!\branch~0_combout  & rfifrdat2_8)

	.dataa(branch),
	.datab(gnd),
	.datac(gnd),
	.datad(rfifrdat2_8),
	.cin(gnd),
	.combout(\RegDat2_ID~8_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~8 .lut_mask = 16'h5500;
defparam \RegDat2_ID~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N1
dffeas \RegDat2_ID[8] (
	.clk(CLK),
	.d(\RegDat2_ID~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[8]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[8] .is_wysiwyg = "true";
defparam \RegDat2_ID[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \Wdata_EX~17 (
// Equation(s):
// \Wdata_EX~17_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_8)) # (!always01 & ((RegDat2_ID[8])))))

	.dataa(Result_EX_8),
	.datab(always0),
	.datac(src2_hazard_t),
	.datad(RegDat2_ID[8]),
	.cin(gnd),
	.combout(\Wdata_EX~17_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~17 .lut_mask = 16'h0B08;
defparam \Wdata_EX~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \Wdata_EX~18 (
// Equation(s):
// \Wdata_EX~18_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~17_combout ) # ((\Equal27~0_combout  & \input_a~111_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(input_a6),
	.datad(\Wdata_EX~17_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~18_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~18 .lut_mask = 16'hAA80;
defparam \Wdata_EX~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \RegDat2_ID~9 (
// Equation(s):
// \RegDat2_ID~9_combout  = (rfifrdat2_9 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_9),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~9_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~9 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N11
dffeas \RegDat2_ID[9] (
	.clk(CLK),
	.d(\RegDat2_ID~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[9]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[9] .is_wysiwyg = "true";
defparam \RegDat2_ID[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \Wdata_EX~19 (
// Equation(s):
// \Wdata_EX~19_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_9))) # (!always01 & (RegDat2_ID[9]))))

	.dataa(src2_hazard_t),
	.datab(RegDat2_ID[9]),
	.datac(Result_EX_9),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~19_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~19 .lut_mask = 16'h5044;
defparam \Wdata_EX~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \Wdata_EX~20 (
// Equation(s):
// \Wdata_EX~20_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~19_combout ) # ((\input_a~108_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(input_a5),
	.datac(Equal27),
	.datad(\Wdata_EX~19_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~20_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~20 .lut_mask = 16'hAA80;
defparam \Wdata_EX~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \RegDat2_ID~10 (
// Equation(s):
// \RegDat2_ID~10_combout  = (!\branch~0_combout  & rfifrdat2_10)

	.dataa(gnd),
	.datab(branch),
	.datac(gnd),
	.datad(rfifrdat2_10),
	.cin(gnd),
	.combout(\RegDat2_ID~10_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~10 .lut_mask = 16'h3300;
defparam \RegDat2_ID~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N29
dffeas \RegDat2_ID[10] (
	.clk(CLK),
	.d(\RegDat2_ID~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[10]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[10] .is_wysiwyg = "true";
defparam \RegDat2_ID[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \Wdata_EX~21 (
// Equation(s):
// \Wdata_EX~21_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_10))) # (!always01 & (RegDat2_ID[10]))))

	.dataa(always0),
	.datab(RegDat2_ID[10]),
	.datac(Result_EX_10),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~21_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~21 .lut_mask = 16'h00E4;
defparam \Wdata_EX~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \Wdata_EX~22 (
// Equation(s):
// \Wdata_EX~22_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~21_combout ) # ((\input_a~105_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~21_combout ),
	.datab(input_a4),
	.datac(\Wdata_EX~0_combout ),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~22_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~22 .lut_mask = 16'hE0A0;
defparam \Wdata_EX~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \RegDat2_ID~11 (
// Equation(s):
// \RegDat2_ID~11_combout  = (rfifrdat2_11 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_11),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~11_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~11 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N29
dffeas \RegDat2_ID[11] (
	.clk(CLK),
	.d(\RegDat2_ID~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[11]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[11] .is_wysiwyg = "true";
defparam \RegDat2_ID[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \Wdata_EX~23 (
// Equation(s):
// \Wdata_EX~23_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_11)) # (!always01 & ((RegDat2_ID[11])))))

	.dataa(always0),
	.datab(src2_hazard_t),
	.datac(Result_EX_11),
	.datad(RegDat2_ID[11]),
	.cin(gnd),
	.combout(\Wdata_EX~23_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~23 .lut_mask = 16'h3120;
defparam \Wdata_EX~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \Wdata_EX~24 (
// Equation(s):
// \Wdata_EX~24_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~23_combout ) # ((\Equal27~0_combout  & \input_a~102_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(\Wdata_EX~23_combout ),
	.datad(input_a3),
	.cin(gnd),
	.combout(\Wdata_EX~24_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~24 .lut_mask = 16'hA8A0;
defparam \Wdata_EX~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \RegDat2_ID~12 (
// Equation(s):
// \RegDat2_ID~12_combout  = (!\branch~0_combout  & rfifrdat2_12)

	.dataa(gnd),
	.datab(branch),
	.datac(gnd),
	.datad(rfifrdat2_12),
	.cin(gnd),
	.combout(\RegDat2_ID~12_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~12 .lut_mask = 16'h3300;
defparam \RegDat2_ID~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N17
dffeas \RegDat2_ID[12] (
	.clk(CLK),
	.d(\RegDat2_ID~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[12]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[12] .is_wysiwyg = "true";
defparam \RegDat2_ID[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \Wdata_EX~25 (
// Equation(s):
// \Wdata_EX~25_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_12)) # (!always01 & ((RegDat2_ID[12])))))

	.dataa(Result_EX_12),
	.datab(src2_hazard_t),
	.datac(RegDat2_ID[12]),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~25_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~25 .lut_mask = 16'h2230;
defparam \Wdata_EX~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \Wdata_EX~26 (
// Equation(s):
// \Wdata_EX~26_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~25_combout ) # ((\input_a~99_combout  & \Equal27~0_combout ))))

	.dataa(input_a2),
	.datab(\Wdata_EX~25_combout ),
	.datac(Equal27),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~26_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~26 .lut_mask = 16'hEC00;
defparam \Wdata_EX~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \Wdata_EX~27 (
// Equation(s):
// \Wdata_EX~27_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_13))) # (!always01 & (RegDat2_ID[13]))))

	.dataa(RegDat2_ID[13]),
	.datab(Result_EX_13),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~27_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~27 .lut_mask = 16'h0C0A;
defparam \Wdata_EX~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \Wdata_EX~28 (
// Equation(s):
// \Wdata_EX~28_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~27_combout ) # ((\Equal27~0_combout  & \input_a~96_combout ))))

	.dataa(\Wdata_EX~27_combout ),
	.datab(Equal27),
	.datac(input_a1),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~28_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~28 .lut_mask = 16'hEA00;
defparam \Wdata_EX~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \RegDat2_ID~14 (
// Equation(s):
// \RegDat2_ID~14_combout  = (!\branch~0_combout  & rfifrdat2_14)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_14),
	.cin(gnd),
	.combout(\RegDat2_ID~14_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~14 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N11
dffeas \RegDat2_ID[14] (
	.clk(CLK),
	.d(\RegDat2_ID~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[14]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[14] .is_wysiwyg = "true";
defparam \RegDat2_ID[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \Wdata_EX~29 (
// Equation(s):
// \Wdata_EX~29_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_14)) # (!always01 & ((RegDat2_ID[14])))))

	.dataa(Result_EX_14),
	.datab(always0),
	.datac(src2_hazard_t),
	.datad(RegDat2_ID[14]),
	.cin(gnd),
	.combout(\Wdata_EX~29_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~29 .lut_mask = 16'h0B08;
defparam \Wdata_EX~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \Wdata_EX~30 (
// Equation(s):
// \Wdata_EX~30_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~29_combout ) # ((\input_b~55_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(input_b16),
	.datac(Equal27),
	.datad(\Wdata_EX~29_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~30_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~30 .lut_mask = 16'hAA80;
defparam \Wdata_EX~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \RegDat2_ID~15 (
// Equation(s):
// \RegDat2_ID~15_combout  = (rfifrdat2_15 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_15),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~15_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~15 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \RegDat2_ID[15] (
	.clk(CLK),
	.d(\RegDat2_ID~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[15]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[15] .is_wysiwyg = "true";
defparam \RegDat2_ID[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \Wdata_EX~31 (
// Equation(s):
// \Wdata_EX~31_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_15))) # (!always01 & (RegDat2_ID[15]))))

	.dataa(always0),
	.datab(src2_hazard_t),
	.datac(RegDat2_ID[15]),
	.datad(Result_EX_15),
	.cin(gnd),
	.combout(\Wdata_EX~31_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~31 .lut_mask = 16'h3210;
defparam \Wdata_EX~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \Wdata_EX~32 (
// Equation(s):
// \Wdata_EX~32_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~31_combout ) # ((\input_b~52_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(\Wdata_EX~31_combout ),
	.datac(input_b15),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~32_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~32 .lut_mask = 16'hA888;
defparam \Wdata_EX~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N12
cycloneive_lcell_comb \RegDat2_ID~16 (
// Equation(s):
// \RegDat2_ID~16_combout  = (rfifrdat2_16 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_16),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~16_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~16 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N13
dffeas \RegDat2_ID[16] (
	.clk(CLK),
	.d(\RegDat2_ID~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[16]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[16] .is_wysiwyg = "true";
defparam \RegDat2_ID[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N2
cycloneive_lcell_comb \Wdata_EX~33 (
// Equation(s):
// \Wdata_EX~33_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_16)) # (!always01 & ((RegDat2_ID[16])))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(Result_EX_16),
	.datad(RegDat2_ID[16]),
	.cin(gnd),
	.combout(\Wdata_EX~33_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~33 .lut_mask = 16'h5140;
defparam \Wdata_EX~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \Wdata_EX~34 (
// Equation(s):
// \Wdata_EX~34_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~33_combout ) # ((\Equal27~0_combout  & \input_b~49_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(\Wdata_EX~33_combout ),
	.datac(Equal27),
	.datad(input_b14),
	.cin(gnd),
	.combout(\Wdata_EX~34_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~34 .lut_mask = 16'hA888;
defparam \Wdata_EX~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \Wdata_EX~35 (
// Equation(s):
// \Wdata_EX~35_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_17))) # (!always01 & (RegDat2_ID[17]))))

	.dataa(RegDat2_ID[17]),
	.datab(src2_hazard_t),
	.datac(Result_EX_17),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~35_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~35 .lut_mask = 16'h3022;
defparam \Wdata_EX~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \Wdata_EX~36 (
// Equation(s):
// \Wdata_EX~36_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~35_combout ) # ((\input_b~46_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~35_combout ),
	.datab(input_b13),
	.datac(Equal27),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~36_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~36 .lut_mask = 16'hEA00;
defparam \Wdata_EX~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N6
cycloneive_lcell_comb \RegDat2_ID~18 (
// Equation(s):
// \RegDat2_ID~18_combout  = (rfifrdat2_18 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(rfifrdat2_18),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~18_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~18 .lut_mask = 16'h00F0;
defparam \RegDat2_ID~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N7
dffeas \RegDat2_ID[18] (
	.clk(CLK),
	.d(\RegDat2_ID~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[18]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[18] .is_wysiwyg = "true";
defparam \RegDat2_ID[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N4
cycloneive_lcell_comb \Wdata_EX~37 (
// Equation(s):
// \Wdata_EX~37_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_18)) # (!always01 & ((RegDat2_ID[18])))))

	.dataa(src2_hazard_t),
	.datab(always0),
	.datac(Result_EX_18),
	.datad(RegDat2_ID[18]),
	.cin(gnd),
	.combout(\Wdata_EX~37_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~37 .lut_mask = 16'h5140;
defparam \Wdata_EX~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \Wdata_EX~38 (
// Equation(s):
// \Wdata_EX~38_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~37_combout ) # ((\Equal27~0_combout  & \input_b~43_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(input_b12),
	.datad(\Wdata_EX~37_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~38_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~38 .lut_mask = 16'hAA80;
defparam \Wdata_EX~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \RegDat2_ID~19 (
// Equation(s):
// \RegDat2_ID~19_combout  = (rfifrdat2_19 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_19),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~19_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~19 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \RegDat2_ID[19] (
	.clk(CLK),
	.d(\RegDat2_ID~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[19]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[19] .is_wysiwyg = "true";
defparam \RegDat2_ID[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \Wdata_EX~39 (
// Equation(s):
// \Wdata_EX~39_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_19)) # (!always01 & ((RegDat2_ID[19])))))

	.dataa(Result_EX_19),
	.datab(src2_hazard_t),
	.datac(RegDat2_ID[19]),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~39_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~39 .lut_mask = 16'h2230;
defparam \Wdata_EX~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \Wdata_EX~40 (
// Equation(s):
// \Wdata_EX~40_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~39_combout ) # ((\Equal27~0_combout  & \input_b~40_combout ))))

	.dataa(Equal27),
	.datab(\Wdata_EX~0_combout ),
	.datac(\Wdata_EX~39_combout ),
	.datad(input_b11),
	.cin(gnd),
	.combout(\Wdata_EX~40_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~40 .lut_mask = 16'hC8C0;
defparam \Wdata_EX~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \RegDat2_ID~20 (
// Equation(s):
// \RegDat2_ID~20_combout  = (rfifrdat2_20 & !\branch~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(rfifrdat2_20),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~20_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~20 .lut_mask = 16'h00F0;
defparam \RegDat2_ID~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N29
dffeas \RegDat2_ID[20] (
	.clk(CLK),
	.d(\RegDat2_ID~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[20]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[20] .is_wysiwyg = "true";
defparam \RegDat2_ID[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \Wdata_EX~41 (
// Equation(s):
// \Wdata_EX~41_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_20))) # (!always01 & (RegDat2_ID[20]))))

	.dataa(always0),
	.datab(RegDat2_ID[20]),
	.datac(Result_EX_20),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~41_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~41 .lut_mask = 16'h00E4;
defparam \Wdata_EX~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \Wdata_EX~42 (
// Equation(s):
// \Wdata_EX~42_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~41_combout ) # ((\input_b~37_combout  & \Equal27~0_combout ))))

	.dataa(input_b10),
	.datab(Equal27),
	.datac(\Wdata_EX~41_combout ),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~42_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~42 .lut_mask = 16'hF800;
defparam \Wdata_EX~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N30
cycloneive_lcell_comb \RegDat2_ID~21 (
// Equation(s):
// \RegDat2_ID~21_combout  = (rfifrdat2_21 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_21),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDat2_ID~21_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~21 .lut_mask = 16'h0C0C;
defparam \RegDat2_ID~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N31
dffeas \RegDat2_ID[21] (
	.clk(CLK),
	.d(\RegDat2_ID~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[21]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[21] .is_wysiwyg = "true";
defparam \RegDat2_ID[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \Wdata_EX~43 (
// Equation(s):
// \Wdata_EX~43_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_21))) # (!always01 & (RegDat2_ID[21]))))

	.dataa(always0),
	.datab(src2_hazard_t),
	.datac(RegDat2_ID[21]),
	.datad(Result_EX_21),
	.cin(gnd),
	.combout(\Wdata_EX~43_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~43 .lut_mask = 16'h3210;
defparam \Wdata_EX~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \Wdata_EX~44 (
// Equation(s):
// \Wdata_EX~44_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~43_combout ) # ((\Equal27~0_combout  & \input_b~34_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(\Wdata_EX~43_combout ),
	.datad(input_b9),
	.cin(gnd),
	.combout(\Wdata_EX~44_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~44 .lut_mask = 16'hA8A0;
defparam \Wdata_EX~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Wdata_EX~45 (
// Equation(s):
// \Wdata_EX~45_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_22))) # (!always01 & (RegDat2_ID[22]))))

	.dataa(RegDat2_ID[22]),
	.datab(Result_EX_22),
	.datac(always0),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~45_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~45 .lut_mask = 16'h00CA;
defparam \Wdata_EX~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \Wdata_EX~46 (
// Equation(s):
// \Wdata_EX~46_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~45_combout ) # ((\Equal27~0_combout  & \input_b~31_combout ))))

	.dataa(\Wdata_EX~45_combout ),
	.datab(Equal27),
	.datac(input_b8),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~46_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~46 .lut_mask = 16'hEA00;
defparam \Wdata_EX~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \RegDat2_ID~23 (
// Equation(s):
// \RegDat2_ID~23_combout  = (rfifrdat2_23 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_23),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDat2_ID~23_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~23 .lut_mask = 16'h0C0C;
defparam \RegDat2_ID~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N19
dffeas \RegDat2_ID[23] (
	.clk(CLK),
	.d(\RegDat2_ID~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[23]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[23] .is_wysiwyg = "true";
defparam \RegDat2_ID[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \Wdata_EX~47 (
// Equation(s):
// \Wdata_EX~47_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_23))) # (!always01 & (RegDat2_ID[23]))))

	.dataa(always0),
	.datab(RegDat2_ID[23]),
	.datac(Result_EX_23),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~47_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~47 .lut_mask = 16'h00E4;
defparam \Wdata_EX~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \Wdata_EX~48 (
// Equation(s):
// \Wdata_EX~48_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~47_combout ) # ((\Equal27~0_combout  & \input_b~28_combout ))))

	.dataa(\Wdata_EX~47_combout ),
	.datab(Equal27),
	.datac(input_b7),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~48_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~48 .lut_mask = 16'hEA00;
defparam \Wdata_EX~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \RegDat2_ID~24 (
// Equation(s):
// \RegDat2_ID~24_combout  = (!\branch~0_combout  & rfifrdat2_24)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_24),
	.cin(gnd),
	.combout(\RegDat2_ID~24_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~24 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N9
dffeas \RegDat2_ID[24] (
	.clk(CLK),
	.d(\RegDat2_ID~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[24]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[24] .is_wysiwyg = "true";
defparam \RegDat2_ID[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \Wdata_EX~49 (
// Equation(s):
// \Wdata_EX~49_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_24)) # (!always01 & ((RegDat2_ID[24])))))

	.dataa(Result_EX_24),
	.datab(always0),
	.datac(RegDat2_ID[24]),
	.datad(src2_hazard_t),
	.cin(gnd),
	.combout(\Wdata_EX~49_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~49 .lut_mask = 16'h00B8;
defparam \Wdata_EX~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \Wdata_EX~50 (
// Equation(s):
// \Wdata_EX~50_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~49_combout ) # ((\Equal27~0_combout  & \input_b~25_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(\Wdata_EX~49_combout ),
	.datad(input_b6),
	.cin(gnd),
	.combout(\Wdata_EX~50_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~50 .lut_mask = 16'hA8A0;
defparam \Wdata_EX~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \RegDat2_ID~25 (
// Equation(s):
// \RegDat2_ID~25_combout  = (rfifrdat2_25 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_25),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~25_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~25 .lut_mask = 16'h00CC;
defparam \RegDat2_ID~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N15
dffeas \RegDat2_ID[25] (
	.clk(CLK),
	.d(\RegDat2_ID~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[25]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[25] .is_wysiwyg = "true";
defparam \RegDat2_ID[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N22
cycloneive_lcell_comb \Wdata_EX~51 (
// Equation(s):
// \Wdata_EX~51_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_25))) # (!always01 & (RegDat2_ID[25]))))

	.dataa(src2_hazard_t),
	.datab(RegDat2_ID[25]),
	.datac(Result_EX_25),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~51_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~51 .lut_mask = 16'h5044;
defparam \Wdata_EX~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N10
cycloneive_lcell_comb \Wdata_EX~52 (
// Equation(s):
// \Wdata_EX~52_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~51_combout ) # ((\Equal27~0_combout  & \input_b~22_combout ))))

	.dataa(Equal27),
	.datab(input_b5),
	.datac(\Wdata_EX~51_combout ),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~52_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~52 .lut_mask = 16'hF800;
defparam \Wdata_EX~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \Wdata_EX~53 (
// Equation(s):
// \Wdata_EX~53_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_26))) # (!always01 & (RegDat2_ID[26]))))

	.dataa(RegDat2_ID[26]),
	.datab(src2_hazard_t),
	.datac(always0),
	.datad(Result_EX_26),
	.cin(gnd),
	.combout(\Wdata_EX~53_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~53 .lut_mask = 16'h3202;
defparam \Wdata_EX~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \Wdata_EX~54 (
// Equation(s):
// \Wdata_EX~54_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~53_combout ) # ((\input_b~19_combout  & \Equal27~0_combout ))))

	.dataa(input_b4),
	.datab(Equal27),
	.datac(\Wdata_EX~53_combout ),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~54_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~54 .lut_mask = 16'hF800;
defparam \Wdata_EX~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \RegDat2_ID~27 (
// Equation(s):
// \RegDat2_ID~27_combout  = (rfifrdat2_27 & !\branch~0_combout )

	.dataa(rfifrdat2_27),
	.datab(gnd),
	.datac(gnd),
	.datad(branch),
	.cin(gnd),
	.combout(\RegDat2_ID~27_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~27 .lut_mask = 16'h00AA;
defparam \RegDat2_ID~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N27
dffeas \RegDat2_ID[27] (
	.clk(CLK),
	.d(\RegDat2_ID~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[27]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[27] .is_wysiwyg = "true";
defparam \RegDat2_ID[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \Wdata_EX~55 (
// Equation(s):
// \Wdata_EX~55_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_27)) # (!always01 & ((RegDat2_ID[27])))))

	.dataa(Result_EX_27),
	.datab(RegDat2_ID[27]),
	.datac(src2_hazard_t),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~55_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~55 .lut_mask = 16'h0A0C;
defparam \Wdata_EX~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \Wdata_EX~56 (
// Equation(s):
// \Wdata_EX~56_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~55_combout ) # ((\Equal27~0_combout  & \input_b~16_combout ))))

	.dataa(\Wdata_EX~55_combout ),
	.datab(Equal27),
	.datac(input_b3),
	.datad(\Wdata_EX~0_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~56_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~56 .lut_mask = 16'hEA00;
defparam \Wdata_EX~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \RegDat2_ID~28 (
// Equation(s):
// \RegDat2_ID~28_combout  = (!\branch~0_combout  & rfifrdat2_28)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_28),
	.cin(gnd),
	.combout(\RegDat2_ID~28_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~28 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N5
dffeas \RegDat2_ID[28] (
	.clk(CLK),
	.d(\RegDat2_ID~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[28]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[28] .is_wysiwyg = "true";
defparam \RegDat2_ID[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \Wdata_EX~57 (
// Equation(s):
// \Wdata_EX~57_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_28))) # (!always01 & (RegDat2_ID[28]))))

	.dataa(always0),
	.datab(src2_hazard_t),
	.datac(RegDat2_ID[28]),
	.datad(Result_EX_28),
	.cin(gnd),
	.combout(\Wdata_EX~57_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~57 .lut_mask = 16'h3210;
defparam \Wdata_EX~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \Wdata_EX~58 (
// Equation(s):
// \Wdata_EX~58_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~57_combout ) # ((\Equal27~0_combout  & \input_b~13_combout ))))

	.dataa(\Wdata_EX~0_combout ),
	.datab(Equal27),
	.datac(\Wdata_EX~57_combout ),
	.datad(input_b2),
	.cin(gnd),
	.combout(\Wdata_EX~58_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~58 .lut_mask = 16'hA8A0;
defparam \Wdata_EX~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \RegDat2_ID~29 (
// Equation(s):
// \RegDat2_ID~29_combout  = (!\branch~0_combout  & rfifrdat2_29)

	.dataa(gnd),
	.datab(gnd),
	.datac(branch),
	.datad(rfifrdat2_29),
	.cin(gnd),
	.combout(\RegDat2_ID~29_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~29 .lut_mask = 16'h0F00;
defparam \RegDat2_ID~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N19
dffeas \RegDat2_ID[29] (
	.clk(CLK),
	.d(\RegDat2_ID~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[29]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[29] .is_wysiwyg = "true";
defparam \RegDat2_ID[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \Wdata_EX~59 (
// Equation(s):
// \Wdata_EX~59_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_29)) # (!always01 & ((RegDat2_ID[29])))))

	.dataa(always0),
	.datab(Result_EX_29),
	.datac(src2_hazard_t),
	.datad(RegDat2_ID[29]),
	.cin(gnd),
	.combout(\Wdata_EX~59_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~59 .lut_mask = 16'h0D08;
defparam \Wdata_EX~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \Wdata_EX~60 (
// Equation(s):
// \Wdata_EX~60_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~59_combout ) # ((\Equal27~0_combout  & \input_b~10_combout ))))

	.dataa(Equal27),
	.datab(input_b1),
	.datac(\Wdata_EX~0_combout ),
	.datad(\Wdata_EX~59_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~60_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~60 .lut_mask = 16'hF080;
defparam \Wdata_EX~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \RegDat2_ID~30 (
// Equation(s):
// \RegDat2_ID~30_combout  = (rfifrdat2_30 & !\branch~0_combout )

	.dataa(gnd),
	.datab(rfifrdat2_30),
	.datac(branch),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDat2_ID~30_combout ),
	.cout());
// synopsys translate_off
defparam \RegDat2_ID~30 .lut_mask = 16'h0C0C;
defparam \RegDat2_ID~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N15
dffeas \RegDat2_ID[30] (
	.clk(CLK),
	.d(\RegDat2_ID~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\care_ID~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(RegDat2_ID[30]),
	.prn(vcc));
// synopsys translate_off
defparam \RegDat2_ID[30] .is_wysiwyg = "true";
defparam \RegDat2_ID[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \Wdata_EX~61 (
// Equation(s):
// \Wdata_EX~61_combout  = (!src2_hazard_t1 & ((always01 & (Result_EX_30)) # (!always01 & ((RegDat2_ID[30])))))

	.dataa(Result_EX_30),
	.datab(src2_hazard_t),
	.datac(always0),
	.datad(RegDat2_ID[30]),
	.cin(gnd),
	.combout(\Wdata_EX~61_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~61 .lut_mask = 16'h2320;
defparam \Wdata_EX~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \Wdata_EX~62 (
// Equation(s):
// \Wdata_EX~62_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~61_combout ) # ((\input_b~7_combout  & \Equal27~0_combout ))))

	.dataa(\Wdata_EX~61_combout ),
	.datab(input_b),
	.datac(\Wdata_EX~0_combout ),
	.datad(Equal27),
	.cin(gnd),
	.combout(\Wdata_EX~62_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~62 .lut_mask = 16'hE0A0;
defparam \Wdata_EX~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \Wdata_EX~63 (
// Equation(s):
// \Wdata_EX~63_combout  = (!src2_hazard_t1 & ((always01 & ((Result_EX_31))) # (!always01 & (RegDat2_ID[31]))))

	.dataa(RegDat2_ID[31]),
	.datab(src2_hazard_t),
	.datac(Result_EX_31),
	.datad(always0),
	.cin(gnd),
	.combout(\Wdata_EX~63_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~63 .lut_mask = 16'h3022;
defparam \Wdata_EX~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \Wdata_EX~64 (
// Equation(s):
// \Wdata_EX~64_combout  = (\Wdata_EX~0_combout  & ((\Wdata_EX~63_combout ) # ((\Equal27~0_combout  & \input_a~56_combout ))))

	.dataa(Equal27),
	.datab(input_a),
	.datac(\Wdata_EX~0_combout ),
	.datad(\Wdata_EX~63_combout ),
	.cin(gnd),
	.combout(\Wdata_EX~64_combout ),
	.cout());
// synopsys translate_off
defparam \Wdata_EX~64 .lut_mask = 16'hF080;
defparam \Wdata_EX~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \Instr_IF~0 (
// Equation(s):
// \Instr_IF~0_combout  = (!always0 & (ramiframload_30 & (!\branch~0_combout  & always1)))

	.dataa(always02),
	.datab(ramiframload_30),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~0_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~0 .lut_mask = 16'h0400;
defparam \Instr_IF~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \Instr_IF~1 (
// Equation(s):
// \Instr_IF~1_combout  = (always1 & (ramiframload_28 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_28),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~1_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~1 .lut_mask = 16'h0008;
defparam \Instr_IF~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \Instr_IF~2 (
// Equation(s):
// \Instr_IF~2_combout  = (always1 & (ramiframload_26 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_26),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~2_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~2 .lut_mask = 16'h0008;
defparam \Instr_IF~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \Instr_IF~3 (
// Equation(s):
// \Instr_IF~3_combout  = (always1 & (ramiframload_27 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_27),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~3_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~3 .lut_mask = 16'h0008;
defparam \Instr_IF~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \Instr_IF~4 (
// Equation(s):
// \Instr_IF~4_combout  = (!always0 & (!\branch~0_combout  & (ramiframload_29 & always1)))

	.dataa(always02),
	.datab(branch),
	.datac(ramiframload_29),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~4_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~4 .lut_mask = 16'h1000;
defparam \Instr_IF~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N24
cycloneive_lcell_comb \Instr_IF~5 (
// Equation(s):
// \Instr_IF~5_combout  = (always1 & (ramiframload_5 & (!\branch~0_combout  & !always0)))

	.dataa(always1),
	.datab(ramiframload_5),
	.datac(branch),
	.datad(always02),
	.cin(gnd),
	.combout(\Instr_IF~5_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~5 .lut_mask = 16'h0008;
defparam \Instr_IF~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N26
cycloneive_lcell_comb \Instr_IF~6 (
// Equation(s):
// \Instr_IF~6_combout  = (ramiframload_4 & (!always0 & (!\branch~0_combout  & always1)))

	.dataa(ramiframload_4),
	.datab(always02),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~6_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~6 .lut_mask = 16'h0200;
defparam \Instr_IF~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \Instr_IF~7 (
// Equation(s):
// \Instr_IF~7_combout  = (always1 & (ramiframload_2 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_2),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~7_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~7 .lut_mask = 16'h0008;
defparam \Instr_IF~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \Instr_IF~8 (
// Equation(s):
// \Instr_IF~8_combout  = (always1 & (!always0 & (ramiframload_3 & !\branch~0_combout )))

	.dataa(always1),
	.datab(always02),
	.datac(ramiframload_3),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~8_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~8 .lut_mask = 16'h0020;
defparam \Instr_IF~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \Instr_IF~9 (
// Equation(s):
// \Instr_IF~9_combout  = (ramiframload_0 & (!always0 & (!\branch~0_combout  & always1)))

	.dataa(ramiframload_0),
	.datab(always02),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~9_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~9 .lut_mask = 16'h0200;
defparam \Instr_IF~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Instr_IF~10 (
// Equation(s):
// \Instr_IF~10_combout  = (!always0 & (ramiframload_1 & (!\branch~0_combout  & always1)))

	.dataa(always02),
	.datab(ramiframload_1),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~10_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~10 .lut_mask = 16'h0400;
defparam \Instr_IF~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \Instr_IF~11 (
// Equation(s):
// \Instr_IF~11_combout  = (ramiframload_31 & (!\branch~0_combout  & (!always0 & always1)))

	.dataa(ramiframload_31),
	.datab(branch),
	.datac(always02),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~11_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~11 .lut_mask = 16'h0200;
defparam \Instr_IF~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \Instr_IF~12 (
// Equation(s):
// \Instr_IF~12_combout  = (always1 & (ramiframload_16 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_16),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~12_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~12 .lut_mask = 16'h0008;
defparam \Instr_IF~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N20
cycloneive_lcell_comb \Instr_IF~13 (
// Equation(s):
// \Instr_IF~13_combout  = (ramiframload_17 & (!always0 & (always1 & !\branch~0_combout )))

	.dataa(ramiframload_17),
	.datab(always02),
	.datac(always1),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~13_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~13 .lut_mask = 16'h0020;
defparam \Instr_IF~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \Instr_IF~14 (
// Equation(s):
// \Instr_IF~14_combout  = (always1 & (ramiframload_18 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_18),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~14_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~14 .lut_mask = 16'h0008;
defparam \Instr_IF~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N30
cycloneive_lcell_comb \Instr_IF~15 (
// Equation(s):
// \Instr_IF~15_combout  = (!\branch~0_combout  & (ramiframload_19 & (always1 & !always0)))

	.dataa(branch),
	.datab(ramiframload_19),
	.datac(always1),
	.datad(always02),
	.cin(gnd),
	.combout(\Instr_IF~15_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~15 .lut_mask = 16'h0040;
defparam \Instr_IF~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \Instr_IF~16 (
// Equation(s):
// \Instr_IF~16_combout  = (ramiframload_20 & (!always0 & (!\branch~0_combout  & always1)))

	.dataa(ramiframload_20),
	.datab(always02),
	.datac(branch),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~16_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~16 .lut_mask = 16'h0200;
defparam \Instr_IF~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \Instr_IF~18 (
// Equation(s):
// \Instr_IF~18_combout  = (ramiframload_21 & (!always0 & (always1 & !\branch~0_combout )))

	.dataa(ramiframload_21),
	.datab(always02),
	.datac(always1),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~18_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~18 .lut_mask = 16'h0020;
defparam \Instr_IF~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \Instr_IF~19 (
// Equation(s):
// \Instr_IF~19_combout  = (ramiframload_22 & (!\branch~0_combout  & (!always0 & always1)))

	.dataa(ramiframload_22),
	.datab(branch),
	.datac(always02),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~19_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~19 .lut_mask = 16'h0200;
defparam \Instr_IF~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \Instr_IF~20 (
// Equation(s):
// \Instr_IF~20_combout  = (always1 & (!always0 & (ramiframload_24 & !\branch~0_combout )))

	.dataa(always1),
	.datab(always02),
	.datac(ramiframload_24),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~20_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~20 .lut_mask = 16'h0020;
defparam \Instr_IF~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Instr_IF~21 (
// Equation(s):
// \Instr_IF~21_combout  = (always1 & (ramiframload_25 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_25),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~21_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~21 .lut_mask = 16'h0008;
defparam \Instr_IF~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \Instr_IF~22 (
// Equation(s):
// \Instr_IF~22_combout  = (ramiframload_23 & (always1 & (!always0 & !\branch~0_combout )))

	.dataa(ramiframload_23),
	.datab(always1),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~22_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~22 .lut_mask = 16'h0008;
defparam \Instr_IF~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N30
cycloneive_lcell_comb \Instr_IF~27 (
// Equation(s):
// \Instr_IF~27_combout  = (!\branch~0_combout  & (ramiframload_10 & (!always0 & always1)))

	.dataa(branch),
	.datab(ramiframload_10),
	.datac(always02),
	.datad(always1),
	.cin(gnd),
	.combout(\Instr_IF~27_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~27 .lut_mask = 16'h0400;
defparam \Instr_IF~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Instr_IF~28 (
// Equation(s):
// \Instr_IF~28_combout  = (!always0 & (ramiframload_9 & (always1 & !\branch~0_combout )))

	.dataa(always02),
	.datab(ramiframload_9),
	.datac(always1),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~28_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~28 .lut_mask = 16'h0040;
defparam \Instr_IF~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \Instr_IF~29 (
// Equation(s):
// \Instr_IF~29_combout  = (always1 & (ramiframload_8 & (!always0 & !\branch~0_combout )))

	.dataa(always1),
	.datab(ramiframload_8),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~29_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~29 .lut_mask = 16'h0008;
defparam \Instr_IF~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \Instr_IF~30 (
// Equation(s):
// \Instr_IF~30_combout  = (ramiframload_7 & (always1 & (!always0 & !\branch~0_combout )))

	.dataa(ramiframload_7),
	.datab(always1),
	.datac(always02),
	.datad(branch),
	.cin(gnd),
	.combout(\Instr_IF~30_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~30 .lut_mask = 16'h0008;
defparam \Instr_IF~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N6
cycloneive_lcell_comb \Instr_IF~31 (
// Equation(s):
// \Instr_IF~31_combout  = (!\branch~0_combout  & (ramiframload_6 & (always1 & !always0)))

	.dataa(branch),
	.datab(ramiframload_6),
	.datac(always1),
	.datad(always02),
	.cin(gnd),
	.combout(\Instr_IF~31_combout ),
	.cout());
// synopsys translate_off
defparam \Instr_IF~31 .lut_mask = 16'h0040;
defparam \Instr_IF~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	input_a,
	RegWen_MEM,
	RegDst_MEM_0,
	RegDst_MEM_1,
	RegDst_MEM_4,
	RegDst_MEM_3,
	RegDst_MEM_2,
	input_b,
	input_b1,
	input_b2,
	input_b3,
	input_b4,
	input_b5,
	input_b6,
	input_b7,
	input_b8,
	input_b9,
	input_b10,
	input_b11,
	input_b12,
	input_b13,
	input_b14,
	input_b15,
	input_b16,
	input_a1,
	input_a2,
	input_a3,
	input_a4,
	input_a5,
	input_a6,
	input_a7,
	input_a8,
	input_a9,
	input_a10,
	input_a11,
	input_a12,
	input_a13,
	input_a14,
	Instr_IF_16,
	Instr_IF_17,
	Instr_IF_18,
	Instr_IF_19,
	Instr_IF_20,
	rfifrdat2_31,
	Instr_IF_21,
	Instr_IF_22,
	Instr_IF_24,
	Instr_IF_25,
	Instr_IF_23,
	rfifrdat1_31,
	rfifrdat1_311,
	WideOr0,
	rfifrdat1_30,
	rfifrdat1_301,
	rfifrdat2_30,
	rfifrdat1_29,
	rfifrdat1_291,
	rfifrdat2_29,
	rfifrdat1_28,
	rfifrdat1_281,
	rfifrdat2_28,
	rfifrdat1_27,
	rfifrdat1_271,
	rfifrdat2_27,
	rfifrdat1_26,
	rfifrdat1_261,
	rfifrdat2_26,
	rfifrdat1_25,
	rfifrdat1_251,
	rfifrdat2_25,
	rfifrdat1_24,
	rfifrdat1_241,
	rfifrdat2_24,
	rfifrdat1_23,
	rfifrdat1_231,
	rfifrdat2_23,
	rfifrdat1_22,
	rfifrdat1_221,
	rfifrdat2_22,
	rfifrdat1_21,
	rfifrdat1_211,
	rfifrdat2_21,
	rfifrdat1_20,
	rfifrdat1_201,
	rfifrdat2_20,
	rfifrdat1_19,
	rfifrdat1_191,
	rfifrdat2_19,
	rfifrdat1_18,
	rfifrdat1_181,
	rfifrdat2_18,
	rfifrdat1_17,
	rfifrdat1_171,
	rfifrdat2_17,
	rfifrdat1_16,
	rfifrdat1_161,
	rfifrdat2_16,
	rfifrdat1_15,
	rfifrdat1_151,
	rfifrdat2_15,
	rfifrdat1_14,
	rfifrdat1_141,
	rfifrdat2_14,
	rfifrdat2_13,
	rfifrdat1_13,
	rfifrdat1_131,
	rfifrdat2_12,
	rfifrdat1_12,
	rfifrdat1_121,
	rfifrdat2_11,
	rfifrdat1_11,
	rfifrdat1_111,
	rfifrdat2_10,
	rfifrdat1_10,
	rfifrdat1_101,
	rfifrdat2_9,
	rfifrdat1_9,
	rfifrdat1_91,
	rfifrdat2_8,
	rfifrdat1_8,
	rfifrdat1_81,
	rfifrdat2_7,
	rfifrdat1_7,
	rfifrdat1_71,
	rfifrdat2_6,
	rfifrdat1_6,
	rfifrdat1_61,
	rfifrdat2_5,
	rfifrdat1_5,
	rfifrdat1_51,
	rfifrdat2_4,
	rfifrdat1_4,
	rfifrdat1_41,
	rfifrdat2_3,
	rfifrdat1_3,
	rfifrdat1_32,
	rfifrdat2_2,
	rfifrdat1_2,
	rfifrdat1_210,
	rfifrdat2_1,
	rfifrdat1_1,
	rfifrdat1_110,
	rfifrdat2_0,
	rfifrdat1_0,
	rfifrdat1_01,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	input_a;
input 	RegWen_MEM;
input 	RegDst_MEM_0;
input 	RegDst_MEM_1;
input 	RegDst_MEM_4;
input 	RegDst_MEM_3;
input 	RegDst_MEM_2;
input 	input_b;
input 	input_b1;
input 	input_b2;
input 	input_b3;
input 	input_b4;
input 	input_b5;
input 	input_b6;
input 	input_b7;
input 	input_b8;
input 	input_b9;
input 	input_b10;
input 	input_b11;
input 	input_b12;
input 	input_b13;
input 	input_b14;
input 	input_b15;
input 	input_b16;
input 	input_a1;
input 	input_a2;
input 	input_a3;
input 	input_a4;
input 	input_a5;
input 	input_a6;
input 	input_a7;
input 	input_a8;
input 	input_a9;
input 	input_a10;
input 	input_a11;
input 	input_a12;
input 	input_a13;
input 	input_a14;
input 	Instr_IF_16;
input 	Instr_IF_17;
input 	Instr_IF_18;
input 	Instr_IF_19;
input 	Instr_IF_20;
output 	rfifrdat2_31;
input 	Instr_IF_21;
input 	Instr_IF_22;
input 	Instr_IF_24;
input 	Instr_IF_25;
input 	Instr_IF_23;
output 	rfifrdat1_31;
output 	rfifrdat1_311;
output 	WideOr0;
output 	rfifrdat1_30;
output 	rfifrdat1_301;
output 	rfifrdat2_30;
output 	rfifrdat1_29;
output 	rfifrdat1_291;
output 	rfifrdat2_29;
output 	rfifrdat1_28;
output 	rfifrdat1_281;
output 	rfifrdat2_28;
output 	rfifrdat1_27;
output 	rfifrdat1_271;
output 	rfifrdat2_27;
output 	rfifrdat1_26;
output 	rfifrdat1_261;
output 	rfifrdat2_26;
output 	rfifrdat1_25;
output 	rfifrdat1_251;
output 	rfifrdat2_25;
output 	rfifrdat1_24;
output 	rfifrdat1_241;
output 	rfifrdat2_24;
output 	rfifrdat1_23;
output 	rfifrdat1_231;
output 	rfifrdat2_23;
output 	rfifrdat1_22;
output 	rfifrdat1_221;
output 	rfifrdat2_22;
output 	rfifrdat1_21;
output 	rfifrdat1_211;
output 	rfifrdat2_21;
output 	rfifrdat1_20;
output 	rfifrdat1_201;
output 	rfifrdat2_20;
output 	rfifrdat1_19;
output 	rfifrdat1_191;
output 	rfifrdat2_19;
output 	rfifrdat1_18;
output 	rfifrdat1_181;
output 	rfifrdat2_18;
output 	rfifrdat1_17;
output 	rfifrdat1_171;
output 	rfifrdat2_17;
output 	rfifrdat1_16;
output 	rfifrdat1_161;
output 	rfifrdat2_16;
output 	rfifrdat1_15;
output 	rfifrdat1_151;
output 	rfifrdat2_15;
output 	rfifrdat1_14;
output 	rfifrdat1_141;
output 	rfifrdat2_14;
output 	rfifrdat2_13;
output 	rfifrdat1_13;
output 	rfifrdat1_131;
output 	rfifrdat2_12;
output 	rfifrdat1_12;
output 	rfifrdat1_121;
output 	rfifrdat2_11;
output 	rfifrdat1_11;
output 	rfifrdat1_111;
output 	rfifrdat2_10;
output 	rfifrdat1_10;
output 	rfifrdat1_101;
output 	rfifrdat2_9;
output 	rfifrdat1_9;
output 	rfifrdat1_91;
output 	rfifrdat2_8;
output 	rfifrdat1_8;
output 	rfifrdat1_81;
output 	rfifrdat2_7;
output 	rfifrdat1_7;
output 	rfifrdat1_71;
output 	rfifrdat2_6;
output 	rfifrdat1_6;
output 	rfifrdat1_61;
output 	rfifrdat2_5;
output 	rfifrdat1_5;
output 	rfifrdat1_51;
output 	rfifrdat2_4;
output 	rfifrdat1_4;
output 	rfifrdat1_41;
output 	rfifrdat2_3;
output 	rfifrdat1_3;
output 	rfifrdat1_32;
output 	rfifrdat2_2;
output 	rfifrdat1_2;
output 	rfifrdat1_210;
output 	rfifrdat2_1;
output 	rfifrdat1_1;
output 	rfifrdat1_110;
output 	rfifrdat2_0;
output 	rfifrdat1_0;
output 	rfifrdat1_01;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \rfif.rdat2[31]~2_combout ;
wire \regs[29][31]~q ;
wire \rfif.rdat2[31]~3_combout ;
wire \regs[20][31]~q ;
wire \rfif.rdat2[31]~7_combout ;
wire \rfif.rdat2[31]~10_combout ;
wire \regs[1][31]~q ;
wire \regs[0][31]~q ;
wire \rfif.rdat2[31]~14_combout ;
wire \rfif.rdat2[31]~15_combout ;
wire \rfif.rdat2[31]~17_combout ;
wire \rfif.rdat1[31]~14_combout ;
wire \regs[19][30]~q ;
wire \regs[12][30]~q ;
wire \rfif.rdat2[30]~28_combout ;
wire \rfif.rdat2[30]~38_combout ;
wire \regs[21][29]~q ;
wire \regs[17][29]~q ;
wire \rfif.rdat1[29]~42_combout ;
wire \regs[28][29]~q ;
wire \regs[3][29]~q ;
wire \regs[12][29]~q ;
wire \rfif.rdat2[29]~44_combout ;
wire \rfif.rdat2[29]~46_combout ;
wire \rfif.rdat2[29]~47_combout ;
wire \rfif.rdat2[29]~56_combout ;
wire \rfif.rdat2[29]~57_combout ;
wire \rfif.rdat2[29]~59_combout ;
wire \rfif.rdat1[28]~72_combout ;
wire \regs[6][27]~q ;
wire \rfif.rdat1[27]~92_combout ;
wire \regs[18][26]~q ;
wire \regs[3][26]~q ;
wire \rfif.rdat2[26]~105_combout ;
wire \rfif.rdat2[26]~107_combout ;
wire \rfif.rdat2[26]~108_combout ;
wire \rfif.rdat2[26]~122_combout ;
wire \rfif.rdat1[25]~122_combout ;
wire \regs[28][25]~q ;
wire \rfif.rdat1[25]~132_combout ;
wire \rfif.rdat2[25]~140_combout ;
wire \rfif.rdat2[25]~141_combout ;
wire \regs[28][24]~q ;
wire \regs[8][24]~q ;
wire \regs[3][24]~q ;
wire \rfif.rdat2[24]~151_combout ;
wire \rfif.rdat2[24]~152_combout ;
wire \rfif.rdat2[24]~154_combout ;
wire \rfif.rdat2[24]~159_combout ;
wire \rfif.rdat2[24]~160_combout ;
wire \regs[28][23]~q ;
wire \regs[4][23]~q ;
wire \rfif.rdat2[23]~168_combout ;
wire \rfif.rdat2[23]~178_combout ;
wire \rfif.rdat2[23]~180_combout ;
wire \rfif.rdat1[22]~184_combout ;
wire \regs[1][22]~q ;
wire \rfif.rdat2[22]~199_combout ;
wire \rfif.rdat2[22]~201_combout ;
wire \rfif.rdat2[22]~206_combout ;
wire \regs[24][21]~q ;
wire \regs[16][21]~q ;
wire \rfif.rdat1[21]~204_combout ;
wire \rfif.rdat1[21]~214_combout ;
wire \rfif.rdat2[21]~214_combout ;
wire \rfif.rdat2[21]~215_combout ;
wire \rfif.rdat2[21]~220_combout ;
wire \rfif.rdat2[21]~222_combout ;
wire \rfif.rdat2[21]~223_combout ;
wire \regs[16][20]~q ;
wire \rfif.rdat2[20]~235_combout ;
wire \rfif.rdat1[19]~242_combout ;
wire \rfif.rdat1[19]~244_combout ;
wire \rfif.rdat1[19]~252_combout ;
wire \regs[2][19]~q ;
wire \regs[1][19]~q ;
wire \rfif.rdat2[19]~269_combout ;
wire \rfif.rdat2[18]~273_combout ;
wire \regs[16][17]~q ;
wire \rfif.rdat1[17]~284_combout ;
wire \rfif.rdat1[17]~292_combout ;
wire \regs[2][17]~q ;
wire \rfif.rdat2[17]~308_combout ;
wire \rfif.rdat2[17]~309_combout ;
wire \regs[22][16]~q ;
wire \regs[18][16]~q ;
wire \rfif.rdat1[16]~302_combout ;
wire \regs[20][16]~q ;
wire \regs[16][16]~q ;
wire \rfif.rdat1[16]~304_combout ;
wire \regs[3][16]~q ;
wire \rfif.rdat2[16]~317_combout ;
wire \rfif.rdat2[16]~318_combout ;
wire \rfif.rdat2[16]~319_combout ;
wire \rfif.rdat2[16]~327_combout ;
wire \rfif.rdat1[15]~332_combout ;
wire \rfif.rdat2[15]~343_combout ;
wire \regs[16][14]~q ;
wire \rfif.rdat1[14]~344_combout ;
wire \rfif.rdat2[14]~357_combout ;
wire \regs[20][13]~q ;
wire \regs[16][13]~q ;
wire \rfif.rdat2[13]~382_combout ;
wire \rfif.rdat2[13]~383_combout ;
wire \regs[4][13]~q ;
wire \rfif.rdat2[13]~390_combout ;
wire \rfif.rdat2[13]~391_combout ;
wire \rfif.rdat1[13]~364_combout ;
wire \regs[19][12]~q ;
wire \rfif.rdat2[12]~406_combout ;
wire \regs[7][12]~q ;
wire \rfif.rdat2[12]~416_combout ;
wire \rfif.rdat1[12]~394_combout ;
wire \regs[16][11]~q ;
wire \rfif.rdat2[11]~424_combout ;
wire \rfif.rdat2[11]~434_combout ;
wire \rfif.rdat2[11]~435_combout ;
wire \regs[1][10]~q ;
wire \regs[0][10]~q ;
wire \rfif.rdat2[10]~455_combout ;
wire \rfif.rdat2[10]~456_combout ;
wire \rfif.rdat1[10]~432_combout ;
wire \rfif.rdat1[10]~434_combout ;
wire \rfif.rdat2[9]~462_combout ;
wire \rfif.rdat2[9]~464_combout ;
wire \regs[20][9]~q ;
wire \regs[9][9]~q ;
wire \regs[8][9]~q ;
wire \rfif.rdat2[9]~472_combout ;
wire \rfif.rdat1[9]~444_combout ;
wire \rfif.rdat1[9]~454_combout ;
wire \rfif.rdat2[8]~485_combout ;
wire \regs[24][8]~q ;
wire \regs[16][8]~q ;
wire \rfif.rdat2[8]~487_combout ;
wire \rfif.rdat2[8]~488_combout ;
wire \rfif.rdat1[8]~464_combout ;
wire \regs[16][7]~q ;
wire \rfif.rdat2[7]~508_combout ;
wire \regs[28][7]~q ;
wire \rfif.rdat2[7]~509_combout ;
wire \regs[24][6]~q ;
wire \regs[16][6]~q ;
wire \rfif.rdat2[6]~529_combout ;
wire \rfif.rdat2[6]~530_combout ;
wire \rfif.rdat2[6]~532_combout ;
wire \rfif.rdat2[6]~542_combout ;
wire \rfif.rdat1[6]~504_combout ;
wire \rfif.rdat1[6]~512_combout ;
wire \rfif.rdat1[6]~514_combout ;
wire \regs[18][5]~q ;
wire \rfif.rdat2[5]~546_combout ;
wire \regs[17][5]~q ;
wire \rfif.rdat2[5]~548_combout ;
wire \rfif.rdat2[5]~549_combout ;
wire \regs[20][5]~q ;
wire \rfif.rdat2[5]~553_combout ;
wire \rfif.rdat1[5]~522_combout ;
wire \rfif.rdat1[5]~524_combout ;
wire \regs[19][4]~q ;
wire \rfif.rdat2[4]~574_combout ;
wire \rfif.rdat2[4]~579_combout ;
wire \rfif.rdat2[4]~580_combout ;
wire \regs[20][3]~q ;
wire \rfif.rdat2[3]~595_combout ;
wire \rfif.rdat2[3]~598_combout ;
wire \regs[4][3]~q ;
wire \rfif.rdat2[3]~600_combout ;
wire \rfif.rdat2[3]~601_combout ;
wire \regs[0][3]~q ;
wire \rfif.rdat2[3]~602_combout ;
wire \rfif.rdat1[3]~562_combout ;
wire \rfif.rdat1[3]~564_combout ;
wire \regs[19][2]~q ;
wire \rfif.rdat2[2]~616_combout ;
wire \rfif.rdat2[1]~630_combout ;
wire \regs[16][1]~q ;
wire \rfif.rdat2[1]~634_combout ;
wire \rfif.rdat2[1]~637_combout ;
wire \rfif.rdat2[0]~653_combout ;
wire \regs[16][0]~q ;
wire \rfif.rdat2[0]~655_combout ;
wire \regs[19][0]~q ;
wire \rfif.rdat2[0]~658_combout ;
wire \rfif.rdat2[0]~661_combout ;
wire \rfif.rdat2[0]~663_combout ;
wire \rfif.rdat2[0]~664_combout ;
wire \regs[20][31]~feeder_combout ;
wire \regs[1][31]~feeder_combout ;
wire \regs[28][29]~feeder_combout ;
wire \regs[3][26]~feeder_combout ;
wire \regs[28][25]~feeder_combout ;
wire \regs[3][24]~feeder_combout ;
wire \regs[28][24]~feeder_combout ;
wire \regs[28][23]~feeder_combout ;
wire \regs[24][21]~feeder_combout ;
wire \regs[1][19]~feeder_combout ;
wire \regs[2][19]~feeder_combout ;
wire \regs[3][16]~feeder_combout ;
wire \regs[7][12]~feeder_combout ;
wire \regs[9][9]~feeder_combout ;
wire \WideOr1~0_combout ;
wire \WideOr1~combout ;
wire \regs[11][31]~feeder_combout ;
wire \Decoder0~18_combout ;
wire \Decoder0~27_combout ;
wire \regs[11][31]~q ;
wire \Decoder0~2_combout ;
wire \Decoder0~24_combout ;
wire \regs[10][31]~q ;
wire \rfif.rdat2[31]~11_combout ;
wire \Decoder0~8_combout ;
wire \Decoder0~28_combout ;
wire \regs[5][31]~q ;
wire \Decoder0~20_combout ;
wire \Decoder0~31_combout ;
wire \regs[7][31]~q ;
wire \Decoder0~0_combout ;
wire \Decoder0~29_combout ;
wire \regs[6][31]~q ;
wire \Decoder0~12_combout ;
wire \Decoder0~30_combout ;
wire \regs[4][31]~q ;
wire \rfif.rdat2[31]~12_combout ;
wire \rfif.rdat2[31]~13_combout ;
wire \rfif.rdat2[31]~16_combout ;
wire \Decoder0~36_combout ;
wire \regs[13][31]~q ;
wire \regs[15][31]~feeder_combout ;
wire \Decoder0~39_combout ;
wire \regs[15][31]~q ;
wire \rfif.rdat2[31]~18_combout ;
wire \rfif.rdat2[31]~19_combout ;
wire \regs[27][31]~feeder_combout ;
wire \Decoder0~19_combout ;
wire \regs[27][31]~q ;
wire \Decoder0~23_combout ;
wire \regs[31][31]~q ;
wire \rfif.rdat2[31]~8_combout ;
wire \Decoder0~5_combout ;
wire \regs[30][31]~q ;
wire \Decoder0~1_combout ;
wire \regs[22][31]~q ;
wire \Decoder0~4_combout ;
wire \regs[18][31]~q ;
wire \Decoder0~3_combout ;
wire \regs[26][31]~q ;
wire \rfif.rdat2[31]~0_combout ;
wire \rfif.rdat2[31]~1_combout ;
wire \Decoder0~14_combout ;
wire \Decoder0~16_combout ;
wire \regs[16][31]~q ;
wire \Decoder0~15_combout ;
wire \regs[24][31]~q ;
wire \rfif.rdat2[31]~4_combout ;
wire \regs[28][31]~feeder_combout ;
wire \Decoder0~17_combout ;
wire \regs[28][31]~q ;
wire \rfif.rdat2[31]~5_combout ;
wire \rfif.rdat2[31]~6_combout ;
wire \rfif.rdat2[31]~9_combout ;
wire \rfif.rdat1[31]~0_combout ;
wire \rfif.rdat1[31]~1_combout ;
wire \regs[23][31]~feeder_combout ;
wire \Decoder0~21_combout ;
wire \regs[23][31]~q ;
wire \regs[19][31]~feeder_combout ;
wire \Decoder0~22_combout ;
wire \regs[19][31]~q ;
wire \rfif.rdat1[31]~7_combout ;
wire \rfif.rdat1[31]~8_combout ;
wire \Decoder0~6_combout ;
wire \Decoder0~7_combout ;
wire \regs[25][31]~q ;
wire \Decoder0~9_combout ;
wire \regs[21][31]~q ;
wire \Decoder0~10_combout ;
wire \regs[17][31]~q ;
wire \rfif.rdat1[31]~2_combout ;
wire \rfif.rdat1[31]~3_combout ;
wire \rfif.rdat1[31]~4_combout ;
wire \rfif.rdat1[31]~5_combout ;
wire \rfif.rdat1[31]~6_combout ;
wire \regs[8][31]~feeder_combout ;
wire \Decoder0~26_combout ;
wire \regs[8][31]~q ;
wire \Decoder0~25_combout ;
wire \regs[9][31]~q ;
wire \rfif.rdat1[31]~10_combout ;
wire \rfif.rdat1[31]~11_combout ;
wire \rfif.rdat1[31]~12_combout ;
wire \rfif.rdat1[31]~13_combout ;
wire \Decoder0~32_combout ;
wire \regs[2][31]~q ;
wire \regs[3][31]~feeder_combout ;
wire \Decoder0~35_combout ;
wire \regs[3][31]~q ;
wire \rfif.rdat1[31]~15_combout ;
wire \rfif.rdat1[31]~16_combout ;
wire \regs[14][31]~feeder_combout ;
wire \Decoder0~37_combout ;
wire \regs[14][31]~q ;
wire \Decoder0~38_combout ;
wire \regs[12][31]~q ;
wire \rfif.rdat1[31]~17_combout ;
wire \rfif.rdat1[31]~18_combout ;
wire \regs[27][30]~feeder_combout ;
wire \regs[27][30]~q ;
wire \rfif.rdat1[30]~27_combout ;
wire \regs[31][30]~feeder_combout ;
wire \regs[31][30]~q ;
wire \regs[23][30]~feeder_combout ;
wire \regs[23][30]~q ;
wire \rfif.rdat1[30]~28_combout ;
wire \regs[16][30]~q ;
wire \regs[20][30]~feeder_combout ;
wire \Decoder0~13_combout ;
wire \regs[20][30]~q ;
wire \rfif.rdat1[30]~24_combout ;
wire \regs[24][30]~q ;
wire \regs[28][30]~feeder_combout ;
wire \regs[28][30]~q ;
wire \rfif.rdat1[30]~25_combout ;
wire \regs[30][30]~q ;
wire \regs[26][30]~q ;
wire \regs[22][30]~q ;
wire \rfif.rdat1[30]~22_combout ;
wire \rfif.rdat1[30]~23_combout ;
wire \rfif.rdat1[30]~26_combout ;
wire \regs[21][30]~q ;
wire \Decoder0~11_combout ;
wire \regs[29][30]~q ;
wire \regs[17][30]~q ;
wire \regs[25][30]~q ;
wire \rfif.rdat1[30]~20_combout ;
wire \rfif.rdat1[30]~21_combout ;
wire \regs[2][30]~q ;
wire \rfif.rdat1[30]~34_combout ;
wire \Decoder0~33_combout ;
wire \regs[1][30]~q ;
wire \regs[3][30]~q ;
wire \rfif.rdat1[30]~35_combout ;
wire \regs[11][30]~q ;
wire \regs[9][30]~q ;
wire \regs[10][30]~q ;
wire \regs[8][30]~q ;
wire \rfif.rdat1[30]~32_combout ;
wire \rfif.rdat1[30]~33_combout ;
wire \rfif.rdat1[30]~36_combout ;
wire \regs[15][30]~q ;
wire \regs[13][30]~q ;
wire \rfif.rdat1[30]~37_combout ;
wire \regs[14][30]~q ;
wire \rfif.rdat1[30]~38_combout ;
wire \regs[5][30]~feeder_combout ;
wire \regs[5][30]~q ;
wire \regs[4][30]~q ;
wire \rfif.rdat1[30]~30_combout ;
wire \regs[7][30]~q ;
wire \regs[6][30]~q ;
wire \rfif.rdat1[30]~31_combout ;
wire \rfif.rdat2[30]~33_combout ;
wire \rfif.rdat2[30]~34_combout ;
wire \Decoder0~34_combout ;
wire \regs[0][30]~q ;
wire \rfif.rdat2[30]~35_combout ;
wire \rfif.rdat2[30]~36_combout ;
wire \rfif.rdat2[30]~37_combout ;
wire \rfif.rdat2[30]~39_combout ;
wire \rfif.rdat2[30]~31_combout ;
wire \rfif.rdat2[30]~32_combout ;
wire \rfif.rdat2[30]~40_combout ;
wire \rfif.rdat2[30]~21_combout ;
wire \rfif.rdat2[30]~22_combout ;
wire \rfif.rdat2[30]~25_combout ;
wire \rfif.rdat2[30]~26_combout ;
wire \regs[18][30]~q ;
wire \rfif.rdat2[30]~23_combout ;
wire \rfif.rdat2[30]~24_combout ;
wire \rfif.rdat2[30]~27_combout ;
wire \rfif.rdat2[30]~29_combout ;
wire \rfif.rdat2[30]~30_combout ;
wire \regs[26][29]~q ;
wire \regs[18][29]~q ;
wire \rfif.rdat1[29]~40_combout ;
wire \regs[30][29]~q ;
wire \regs[22][29]~q ;
wire \rfif.rdat1[29]~41_combout ;
wire \regs[25][29]~q ;
wire \regs[29][29]~q ;
wire \rfif.rdat1[29]~43_combout ;
wire \regs[24][29]~q ;
wire \regs[16][29]~q ;
wire \rfif.rdat1[29]~44_combout ;
wire \regs[20][29]~feeder_combout ;
wire \regs[20][29]~q ;
wire \rfif.rdat1[29]~45_combout ;
wire \rfif.rdat1[29]~46_combout ;
wire \regs[31][29]~feeder_combout ;
wire \regs[31][29]~q ;
wire \regs[23][29]~feeder_combout ;
wire \regs[23][29]~q ;
wire \regs[19][29]~feeder_combout ;
wire \regs[19][29]~q ;
wire \rfif.rdat1[29]~47_combout ;
wire \regs[27][29]~feeder_combout ;
wire \regs[27][29]~q ;
wire \rfif.rdat1[29]~48_combout ;
wire \regs[14][29]~feeder_combout ;
wire \regs[14][29]~q ;
wire \rfif.rdat1[29]~57_combout ;
wire \regs[15][29]~q ;
wire \regs[13][29]~q ;
wire \rfif.rdat1[29]~58_combout ;
wire \regs[6][29]~feeder_combout ;
wire \regs[6][29]~q ;
wire \rfif.rdat1[29]~52_combout ;
wire \regs[5][29]~q ;
wire \regs[7][29]~q ;
wire \rfif.rdat1[29]~53_combout ;
wire \regs[2][29]~q ;
wire \regs[1][29]~feeder_combout ;
wire \regs[1][29]~q ;
wire \regs[0][29]~q ;
wire \rfif.rdat1[29]~54_combout ;
wire \rfif.rdat1[29]~55_combout ;
wire \rfif.rdat1[29]~56_combout ;
wire \regs[8][29]~feeder_combout ;
wire \regs[8][29]~q ;
wire \regs[9][29]~q ;
wire \rfif.rdat1[29]~50_combout ;
wire \regs[11][29]~q ;
wire \regs[10][29]~feeder_combout ;
wire \regs[10][29]~q ;
wire \rfif.rdat1[29]~51_combout ;
wire \rfif.rdat2[29]~52_combout ;
wire \rfif.rdat2[29]~53_combout ;
wire \regs[4][29]~q ;
wire \rfif.rdat2[29]~54_combout ;
wire \rfif.rdat2[29]~55_combout ;
wire \rfif.rdat2[29]~58_combout ;
wire \rfif.rdat2[29]~60_combout ;
wire \rfif.rdat2[29]~61_combout ;
wire \rfif.rdat2[29]~42_combout ;
wire \rfif.rdat2[29]~43_combout ;
wire \rfif.rdat2[29]~49_combout ;
wire \rfif.rdat2[29]~50_combout ;
wire \rfif.rdat2[29]~45_combout ;
wire \rfif.rdat2[29]~48_combout ;
wire \rfif.rdat2[29]~51_combout ;
wire \regs[24][28]~feeder_combout ;
wire \regs[24][28]~q ;
wire \regs[28][28]~q ;
wire \regs[20][28]~feeder_combout ;
wire \regs[20][28]~q ;
wire \regs[16][28]~q ;
wire \rfif.rdat1[28]~64_combout ;
wire \rfif.rdat1[28]~65_combout ;
wire \regs[22][28]~q ;
wire \rfif.rdat1[28]~62_combout ;
wire \regs[26][28]~q ;
wire \regs[30][28]~q ;
wire \rfif.rdat1[28]~63_combout ;
wire \rfif.rdat1[28]~66_combout ;
wire \regs[31][28]~feeder_combout ;
wire \regs[31][28]~q ;
wire \regs[23][28]~feeder_combout ;
wire \regs[23][28]~q ;
wire \regs[27][28]~feeder_combout ;
wire \regs[27][28]~q ;
wire \regs[19][28]~q ;
wire \rfif.rdat1[28]~67_combout ;
wire \rfif.rdat1[28]~68_combout ;
wire \regs[29][28]~feeder_combout ;
wire \regs[29][28]~q ;
wire \regs[17][28]~feeder_combout ;
wire \regs[17][28]~q ;
wire \regs[25][28]~q ;
wire \rfif.rdat1[28]~60_combout ;
wire \regs[21][28]~q ;
wire \rfif.rdat1[28]~61_combout ;
wire \regs[15][28]~q ;
wire \regs[14][28]~q ;
wire \regs[13][28]~q ;
wire \rfif.rdat1[28]~77_combout ;
wire \rfif.rdat1[28]~78_combout ;
wire \regs[9][28]~q ;
wire \regs[11][28]~q ;
wire \rfif.rdat1[28]~73_combout ;
wire \regs[2][28]~feeder_combout ;
wire \regs[2][28]~q ;
wire \regs[0][28]~q ;
wire \rfif.rdat1[28]~74_combout ;
wire \regs[1][28]~q ;
wire \regs[3][28]~q ;
wire \rfif.rdat1[28]~75_combout ;
wire \rfif.rdat1[28]~76_combout ;
wire \regs[4][28]~q ;
wire \regs[5][28]~q ;
wire \rfif.rdat1[28]~70_combout ;
wire \regs[7][28]~q ;
wire \regs[6][28]~q ;
wire \rfif.rdat1[28]~71_combout ;
wire \regs[12][28]~q ;
wire \rfif.rdat2[28]~80_combout ;
wire \rfif.rdat2[28]~81_combout ;
wire \rfif.rdat2[28]~73_combout ;
wire \rfif.rdat2[28]~74_combout ;
wire \rfif.rdat2[28]~77_combout ;
wire \rfif.rdat2[28]~78_combout ;
wire \regs[8][28]~q ;
wire \regs[10][28]~q ;
wire \rfif.rdat2[28]~75_combout ;
wire \rfif.rdat2[28]~76_combout ;
wire \rfif.rdat2[28]~79_combout ;
wire \rfif.rdat2[28]~82_combout ;
wire \rfif.rdat2[28]~70_combout ;
wire \rfif.rdat2[28]~71_combout ;
wire \rfif.rdat2[28]~63_combout ;
wire \rfif.rdat2[28]~64_combout ;
wire \rfif.rdat2[28]~67_combout ;
wire \rfif.rdat2[28]~68_combout ;
wire \regs[18][28]~q ;
wire \rfif.rdat2[28]~65_combout ;
wire \rfif.rdat2[28]~66_combout ;
wire \rfif.rdat2[28]~69_combout ;
wire \rfif.rdat2[28]~72_combout ;
wire \regs[23][27]~feeder_combout ;
wire \regs[23][27]~q ;
wire \regs[19][27]~q ;
wire \rfif.rdat1[27]~87_combout ;
wire \regs[31][27]~q ;
wire \regs[27][27]~q ;
wire \rfif.rdat1[27]~88_combout ;
wire \regs[22][27]~q ;
wire \regs[30][27]~q ;
wire \regs[18][27]~q ;
wire \regs[26][27]~q ;
wire \rfif.rdat1[27]~80_combout ;
wire \rfif.rdat1[27]~81_combout ;
wire \regs[20][27]~feeder_combout ;
wire \regs[20][27]~q ;
wire \regs[16][27]~q ;
wire \regs[24][27]~q ;
wire \rfif.rdat1[27]~84_combout ;
wire \rfif.rdat1[27]~85_combout ;
wire \regs[25][27]~q ;
wire \regs[17][27]~q ;
wire \regs[21][27]~q ;
wire \rfif.rdat1[27]~82_combout ;
wire \rfif.rdat1[27]~83_combout ;
wire \rfif.rdat1[27]~86_combout ;
wire \regs[1][27]~feeder_combout ;
wire \regs[1][27]~q ;
wire \regs[0][27]~q ;
wire \rfif.rdat1[27]~94_combout ;
wire \regs[2][27]~q ;
wire \regs[3][27]~q ;
wire \rfif.rdat1[27]~95_combout ;
wire \regs[5][27]~q ;
wire \regs[7][27]~q ;
wire \rfif.rdat1[27]~93_combout ;
wire \rfif.rdat1[27]~96_combout ;
wire \regs[15][27]~feeder_combout ;
wire \regs[15][27]~q ;
wire \regs[13][27]~q ;
wire \regs[14][27]~feeder_combout ;
wire \regs[14][27]~q ;
wire \regs[12][27]~q ;
wire \rfif.rdat1[27]~97_combout ;
wire \rfif.rdat1[27]~98_combout ;
wire \regs[11][27]~feeder_combout ;
wire \regs[11][27]~q ;
wire \regs[10][27]~feeder_combout ;
wire \regs[10][27]~q ;
wire \regs[9][27]~q ;
wire \regs[8][27]~q ;
wire \rfif.rdat1[27]~90_combout ;
wire \rfif.rdat1[27]~91_combout ;
wire \rfif.rdat2[27]~94_combout ;
wire \rfif.rdat2[27]~95_combout ;
wire \rfif.rdat2[27]~101_combout ;
wire \rfif.rdat2[27]~102_combout ;
wire \regs[4][27]~q ;
wire \rfif.rdat2[27]~96_combout ;
wire \rfif.rdat2[27]~97_combout ;
wire \rfif.rdat2[27]~98_combout ;
wire \rfif.rdat2[27]~99_combout ;
wire \rfif.rdat2[27]~100_combout ;
wire \rfif.rdat2[27]~103_combout ;
wire \rfif.rdat2[27]~91_combout ;
wire \rfif.rdat2[27]~92_combout ;
wire \rfif.rdat2[27]~84_combout ;
wire \rfif.rdat2[27]~85_combout ;
wire \regs[29][27]~q ;
wire \rfif.rdat2[27]~86_combout ;
wire \rfif.rdat2[27]~87_combout ;
wire \regs[28][27]~feeder_combout ;
wire \regs[28][27]~q ;
wire \rfif.rdat2[27]~88_combout ;
wire \rfif.rdat2[27]~89_combout ;
wire \rfif.rdat2[27]~90_combout ;
wire \rfif.rdat2[27]~93_combout ;
wire \regs[31][26]~q ;
wire \regs[23][26]~q ;
wire \regs[19][26]~q ;
wire \regs[27][26]~feeder_combout ;
wire \regs[27][26]~q ;
wire \rfif.rdat1[26]~107_combout ;
wire \rfif.rdat1[26]~108_combout ;
wire \regs[21][26]~q ;
wire \regs[17][26]~q ;
wire \regs[25][26]~q ;
wire \rfif.rdat1[26]~100_combout ;
wire \regs[29][26]~q ;
wire \rfif.rdat1[26]~101_combout ;
wire \regs[16][26]~q ;
wire \regs[20][26]~q ;
wire \rfif.rdat1[26]~104_combout ;
wire \regs[24][26]~q ;
wire \regs[28][26]~q ;
wire \rfif.rdat1[26]~105_combout ;
wire \regs[30][26]~q ;
wire \regs[26][26]~q ;
wire \regs[22][26]~q ;
wire \rfif.rdat1[26]~102_combout ;
wire \rfif.rdat1[26]~103_combout ;
wire \rfif.rdat1[26]~106_combout ;
wire \regs[6][26]~q ;
wire \regs[7][26]~q ;
wire \regs[5][26]~q ;
wire \rfif.rdat1[26]~110_combout ;
wire \rfif.rdat1[26]~111_combout ;
wire \regs[14][26]~feeder_combout ;
wire \regs[14][26]~q ;
wire \regs[15][26]~q ;
wire \regs[12][26]~q ;
wire \regs[13][26]~q ;
wire \rfif.rdat1[26]~117_combout ;
wire \rfif.rdat1[26]~118_combout ;
wire \regs[0][26]~q ;
wire \regs[2][26]~q ;
wire \rfif.rdat1[26]~114_combout ;
wire \regs[1][26]~feeder_combout ;
wire \regs[1][26]~q ;
wire \rfif.rdat1[26]~115_combout ;
wire \regs[11][26]~q ;
wire \regs[10][26]~q ;
wire \regs[8][26]~q ;
wire \rfif.rdat1[26]~112_combout ;
wire \regs[9][26]~feeder_combout ;
wire \regs[9][26]~q ;
wire \rfif.rdat1[26]~113_combout ;
wire \rfif.rdat1[26]~116_combout ;
wire \regs[4][26]~q ;
wire \rfif.rdat2[26]~115_combout ;
wire \rfif.rdat2[26]~116_combout ;
wire \rfif.rdat2[26]~123_combout ;
wire \rfif.rdat2[26]~117_combout ;
wire \rfif.rdat2[26]~118_combout ;
wire \rfif.rdat2[26]~119_combout ;
wire \rfif.rdat2[26]~120_combout ;
wire \rfif.rdat2[26]~121_combout ;
wire \rfif.rdat2[26]~124_combout ;
wire \rfif.rdat2[26]~106_combout ;
wire \rfif.rdat2[26]~109_combout ;
wire \rfif.rdat2[26]~110_combout ;
wire \rfif.rdat2[26]~111_combout ;
wire \rfif.rdat2[26]~112_combout ;
wire \rfif.rdat2[26]~113_combout ;
wire \rfif.rdat2[26]~114_combout ;
wire \regs[23][25]~q ;
wire \regs[19][25]~q ;
wire \rfif.rdat1[25]~127_combout ;
wire \regs[27][25]~q ;
wire \regs[31][25]~q ;
wire \rfif.rdat1[25]~128_combout ;
wire \regs[26][25]~q ;
wire \regs[18][25]~q ;
wire \rfif.rdat1[25]~120_combout ;
wire \regs[30][25]~q ;
wire \regs[22][25]~q ;
wire \rfif.rdat1[25]~121_combout ;
wire \regs[29][25]~q ;
wire \regs[25][25]~q ;
wire \rfif.rdat1[25]~123_combout ;
wire \regs[20][25]~feeder_combout ;
wire \regs[20][25]~q ;
wire \regs[16][25]~q ;
wire \regs[24][25]~q ;
wire \rfif.rdat1[25]~124_combout ;
wire \rfif.rdat1[25]~125_combout ;
wire \rfif.rdat1[25]~126_combout ;
wire \regs[3][25]~feeder_combout ;
wire \regs[3][25]~q ;
wire \regs[2][25]~q ;
wire \regs[1][25]~q ;
wire \regs[0][25]~q ;
wire \rfif.rdat1[25]~134_combout ;
wire \rfif.rdat1[25]~135_combout ;
wire \regs[7][25]~feeder_combout ;
wire \regs[7][25]~q ;
wire \regs[5][25]~q ;
wire \rfif.rdat1[25]~133_combout ;
wire \rfif.rdat1[25]~136_combout ;
wire \regs[8][25]~q ;
wire \regs[9][25]~feeder_combout ;
wire \regs[9][25]~q ;
wire \rfif.rdat1[25]~130_combout ;
wire \regs[10][25]~q ;
wire \regs[11][25]~feeder_combout ;
wire \regs[11][25]~q ;
wire \rfif.rdat1[25]~131_combout ;
wire \regs[15][25]~feeder_combout ;
wire \regs[15][25]~q ;
wire \regs[12][25]~q ;
wire \regs[14][25]~q ;
wire \rfif.rdat1[25]~137_combout ;
wire \regs[13][25]~q ;
wire \rfif.rdat1[25]~138_combout ;
wire \rfif.rdat2[25]~136_combout ;
wire \rfif.rdat2[25]~137_combout ;
wire \rfif.rdat2[25]~143_combout ;
wire \rfif.rdat2[25]~144_combout ;
wire \regs[4][25]~q ;
wire \regs[6][25]~q ;
wire \rfif.rdat2[25]~138_combout ;
wire \rfif.rdat2[25]~139_combout ;
wire \rfif.rdat2[25]~142_combout ;
wire \rfif.rdat2[25]~145_combout ;
wire \rfif.rdat2[25]~126_combout ;
wire \rfif.rdat2[25]~127_combout ;
wire \rfif.rdat2[25]~133_combout ;
wire \rfif.rdat2[25]~134_combout ;
wire \regs[17][25]~q ;
wire \regs[21][25]~q ;
wire \rfif.rdat2[25]~128_combout ;
wire \rfif.rdat2[25]~129_combout ;
wire \rfif.rdat2[25]~130_combout ;
wire \rfif.rdat2[25]~131_combout ;
wire \rfif.rdat2[25]~132_combout ;
wire \rfif.rdat2[25]~135_combout ;
wire \regs[21][24]~q ;
wire \regs[17][24]~q ;
wire \regs[25][24]~q ;
wire \rfif.rdat1[24]~140_combout ;
wire \regs[29][24]~q ;
wire \rfif.rdat1[24]~141_combout ;
wire \regs[24][24]~feeder_combout ;
wire \regs[24][24]~q ;
wire \regs[20][24]~q ;
wire \regs[16][24]~q ;
wire \rfif.rdat1[24]~144_combout ;
wire \rfif.rdat1[24]~145_combout ;
wire \regs[26][24]~q ;
wire \regs[22][24]~q ;
wire \rfif.rdat1[24]~142_combout ;
wire \rfif.rdat1[24]~143_combout ;
wire \rfif.rdat1[24]~146_combout ;
wire \regs[23][24]~feeder_combout ;
wire \regs[23][24]~q ;
wire \regs[27][24]~feeder_combout ;
wire \regs[27][24]~q ;
wire \regs[19][24]~q ;
wire \rfif.rdat1[24]~147_combout ;
wire \regs[31][24]~feeder_combout ;
wire \regs[31][24]~q ;
wire \rfif.rdat1[24]~148_combout ;
wire \regs[15][24]~feeder_combout ;
wire \regs[15][24]~q ;
wire \regs[12][24]~q ;
wire \regs[13][24]~q ;
wire \rfif.rdat1[24]~157_combout ;
wire \regs[14][24]~feeder_combout ;
wire \regs[14][24]~q ;
wire \rfif.rdat1[24]~158_combout ;
wire \regs[6][24]~q ;
wire \regs[7][24]~q ;
wire \regs[5][24]~q ;
wire \rfif.rdat1[24]~150_combout ;
wire \rfif.rdat1[24]~151_combout ;
wire \regs[1][24]~feeder_combout ;
wire \regs[1][24]~q ;
wire \regs[2][24]~q ;
wire \regs[0][24]~q ;
wire \rfif.rdat1[24]~154_combout ;
wire \rfif.rdat1[24]~155_combout ;
wire \regs[11][24]~q ;
wire \regs[9][24]~q ;
wire \regs[10][24]~feeder_combout ;
wire \regs[10][24]~q ;
wire \rfif.rdat1[24]~152_combout ;
wire \rfif.rdat1[24]~153_combout ;
wire \rfif.rdat1[24]~156_combout ;
wire \rfif.rdat2[24]~147_combout ;
wire \rfif.rdat2[24]~148_combout ;
wire \rfif.rdat2[24]~155_combout ;
wire \regs[30][24]~q ;
wire \regs[18][24]~q ;
wire \rfif.rdat2[24]~149_combout ;
wire \rfif.rdat2[24]~150_combout ;
wire \rfif.rdat2[24]~153_combout ;
wire \rfif.rdat2[24]~156_combout ;
wire \rfif.rdat2[24]~164_combout ;
wire \rfif.rdat2[24]~165_combout ;
wire \rfif.rdat2[24]~161_combout ;
wire \rfif.rdat2[24]~162_combout ;
wire \rfif.rdat2[24]~163_combout ;
wire \regs[4][24]~q ;
wire \rfif.rdat2[24]~157_combout ;
wire \rfif.rdat2[24]~158_combout ;
wire \rfif.rdat2[24]~166_combout ;
wire \regs[26][23]~q ;
wire \regs[18][23]~q ;
wire \rfif.rdat1[23]~160_combout ;
wire \regs[22][23]~q ;
wire \regs[30][23]~q ;
wire \rfif.rdat1[23]~161_combout ;
wire \regs[19][23]~q ;
wire \regs[23][23]~feeder_combout ;
wire \regs[23][23]~q ;
wire \rfif.rdat1[23]~167_combout ;
wire \regs[31][23]~q ;
wire \regs[27][23]~q ;
wire \rfif.rdat1[23]~168_combout ;
wire \regs[25][23]~q ;
wire \regs[21][23]~q ;
wire \regs[17][23]~q ;
wire \rfif.rdat1[23]~162_combout ;
wire \rfif.rdat1[23]~163_combout ;
wire \regs[20][23]~q ;
wire \regs[24][23]~feeder_combout ;
wire \regs[24][23]~q ;
wire \regs[16][23]~q ;
wire \rfif.rdat1[23]~164_combout ;
wire \rfif.rdat1[23]~165_combout ;
wire \rfif.rdat1[23]~166_combout ;
wire \regs[0][23]~q ;
wire \regs[1][23]~feeder_combout ;
wire \regs[1][23]~q ;
wire \rfif.rdat1[23]~174_combout ;
wire \regs[3][23]~q ;
wire \regs[2][23]~q ;
wire \rfif.rdat1[23]~175_combout ;
wire \regs[5][23]~q ;
wire \regs[6][23]~q ;
wire \rfif.rdat1[23]~172_combout ;
wire \rfif.rdat1[23]~173_combout ;
wire \rfif.rdat1[23]~176_combout ;
wire \regs[14][23]~q ;
wire \regs[12][23]~q ;
wire \rfif.rdat1[23]~177_combout ;
wire \regs[15][23]~q ;
wire \regs[13][23]~q ;
wire \rfif.rdat1[23]~178_combout ;
wire \regs[10][23]~q ;
wire \regs[9][23]~q ;
wire \regs[8][23]~q ;
wire \rfif.rdat1[23]~170_combout ;
wire \regs[11][23]~q ;
wire \rfif.rdat1[23]~171_combout ;
wire \rfif.rdat2[23]~179_combout ;
wire \rfif.rdat2[23]~185_combout ;
wire \rfif.rdat2[23]~186_combout ;
wire \rfif.rdat2[23]~182_combout ;
wire \rfif.rdat2[23]~183_combout ;
wire \regs[7][23]~q ;
wire \rfif.rdat2[23]~181_combout ;
wire \rfif.rdat2[23]~184_combout ;
wire \rfif.rdat2[23]~187_combout ;
wire \rfif.rdat2[23]~169_combout ;
wire \rfif.rdat2[23]~175_combout ;
wire \rfif.rdat2[23]~176_combout ;
wire \regs[29][23]~q ;
wire \rfif.rdat2[23]~170_combout ;
wire \rfif.rdat2[23]~171_combout ;
wire \rfif.rdat2[23]~172_combout ;
wire \rfif.rdat2[23]~173_combout ;
wire \rfif.rdat2[23]~174_combout ;
wire \rfif.rdat2[23]~177_combout ;
wire \regs[24][22]~feeder_combout ;
wire \regs[24][22]~q ;
wire \regs[28][22]~feeder_combout ;
wire \regs[28][22]~q ;
wire \rfif.rdat1[22]~185_combout ;
wire \regs[22][22]~q ;
wire \regs[18][22]~q ;
wire \rfif.rdat1[22]~182_combout ;
wire \regs[26][22]~q ;
wire \rfif.rdat1[22]~183_combout ;
wire \rfif.rdat1[22]~186_combout ;
wire \regs[17][22]~q ;
wire \regs[25][22]~q ;
wire \rfif.rdat1[22]~180_combout ;
wire \regs[29][22]~q ;
wire \regs[21][22]~q ;
wire \rfif.rdat1[22]~181_combout ;
wire \regs[23][22]~feeder_combout ;
wire \regs[23][22]~q ;
wire \regs[31][22]~q ;
wire \regs[27][22]~q ;
wire \regs[19][22]~q ;
wire \rfif.rdat1[22]~187_combout ;
wire \rfif.rdat1[22]~188_combout ;
wire \regs[14][22]~feeder_combout ;
wire \regs[14][22]~q ;
wire \regs[12][22]~q ;
wire \regs[13][22]~q ;
wire \rfif.rdat1[22]~197_combout ;
wire \regs[15][22]~q ;
wire \rfif.rdat1[22]~198_combout ;
wire \regs[3][22]~feeder_combout ;
wire \regs[3][22]~q ;
wire \regs[2][22]~q ;
wire \regs[0][22]~q ;
wire \rfif.rdat1[22]~194_combout ;
wire \rfif.rdat1[22]~195_combout ;
wire \regs[10][22]~q ;
wire \regs[8][22]~q ;
wire \rfif.rdat1[22]~192_combout ;
wire \regs[9][22]~q ;
wire \rfif.rdat1[22]~193_combout ;
wire \rfif.rdat1[22]~196_combout ;
wire \regs[6][22]~q ;
wire \regs[7][22]~q ;
wire \regs[5][22]~q ;
wire \regs[4][22]~q ;
wire \rfif.rdat1[22]~190_combout ;
wire \rfif.rdat1[22]~191_combout ;
wire \rfif.rdat2[22]~189_combout ;
wire \rfif.rdat2[22]~190_combout ;
wire \rfif.rdat2[22]~196_combout ;
wire \rfif.rdat2[22]~197_combout ;
wire \regs[16][22]~q ;
wire \regs[20][22]~q ;
wire \rfif.rdat2[22]~193_combout ;
wire \rfif.rdat2[22]~194_combout ;
wire \regs[30][22]~q ;
wire \rfif.rdat2[22]~191_combout ;
wire \rfif.rdat2[22]~192_combout ;
wire \rfif.rdat2[22]~195_combout ;
wire \rfif.rdat2[22]~198_combout ;
wire \regs[11][22]~q ;
wire \rfif.rdat2[22]~202_combout ;
wire \rfif.rdat2[22]~203_combout ;
wire \rfif.rdat2[22]~204_combout ;
wire \rfif.rdat2[22]~205_combout ;
wire \rfif.rdat2[22]~200_combout ;
wire \rfif.rdat2[22]~207_combout ;
wire \rfif.rdat2[22]~208_combout ;
wire \regs[20][21]~q ;
wire \regs[28][21]~feeder_combout ;
wire \regs[28][21]~q ;
wire \rfif.rdat1[21]~205_combout ;
wire \regs[25][21]~q ;
wire \regs[21][21]~q ;
wire \rfif.rdat1[21]~202_combout ;
wire \rfif.rdat1[21]~203_combout ;
wire \rfif.rdat1[21]~206_combout ;
wire \regs[27][21]~feeder_combout ;
wire \regs[27][21]~q ;
wire \regs[19][21]~q ;
wire \regs[23][21]~q ;
wire \rfif.rdat1[21]~207_combout ;
wire \regs[31][21]~q ;
wire \rfif.rdat1[21]~208_combout ;
wire \regs[22][21]~q ;
wire \regs[30][21]~q ;
wire \regs[26][21]~q ;
wire \regs[18][21]~q ;
wire \rfif.rdat1[21]~200_combout ;
wire \rfif.rdat1[21]~201_combout ;
wire \regs[7][21]~feeder_combout ;
wire \regs[7][21]~q ;
wire \regs[6][21]~q ;
wire \regs[4][21]~q ;
wire \rfif.rdat1[21]~212_combout ;
wire \regs[5][21]~feeder_combout ;
wire \regs[5][21]~q ;
wire \rfif.rdat1[21]~213_combout ;
wire \regs[3][21]~feeder_combout ;
wire \regs[3][21]~q ;
wire \regs[2][21]~q ;
wire \rfif.rdat1[21]~215_combout ;
wire \rfif.rdat1[21]~216_combout ;
wire \regs[8][21]~q ;
wire \regs[9][21]~q ;
wire \rfif.rdat1[21]~210_combout ;
wire \regs[11][21]~q ;
wire \regs[10][21]~q ;
wire \rfif.rdat1[21]~211_combout ;
wire \regs[15][21]~q ;
wire \regs[14][21]~q ;
wire \regs[12][21]~q ;
wire \rfif.rdat1[21]~217_combout ;
wire \regs[13][21]~q ;
wire \rfif.rdat1[21]~218_combout ;
wire \rfif.rdat2[21]~227_combout ;
wire \rfif.rdat2[21]~228_combout ;
wire \rfif.rdat2[21]~221_combout ;
wire \regs[1][21]~feeder_combout ;
wire \regs[1][21]~q ;
wire \regs[0][21]~q ;
wire \rfif.rdat2[21]~224_combout ;
wire \rfif.rdat2[21]~225_combout ;
wire \rfif.rdat2[21]~226_combout ;
wire \rfif.rdat2[21]~229_combout ;
wire \rfif.rdat2[21]~217_combout ;
wire \rfif.rdat2[21]~218_combout ;
wire \rfif.rdat2[21]~210_combout ;
wire \rfif.rdat2[21]~211_combout ;
wire \regs[29][21]~q ;
wire \regs[17][21]~q ;
wire \rfif.rdat2[21]~212_combout ;
wire \rfif.rdat2[21]~213_combout ;
wire \rfif.rdat2[21]~216_combout ;
wire \rfif.rdat2[21]~219_combout ;
wire \regs[27][20]~q ;
wire \regs[19][20]~q ;
wire \rfif.rdat1[20]~227_combout ;
wire \regs[23][20]~q ;
wire \regs[31][20]~q ;
wire \rfif.rdat1[20]~228_combout ;
wire \regs[21][20]~q ;
wire \regs[29][20]~q ;
wire \regs[17][20]~q ;
wire \regs[25][20]~q ;
wire \rfif.rdat1[20]~220_combout ;
wire \rfif.rdat1[20]~221_combout ;
wire \regs[24][20]~feeder_combout ;
wire \regs[24][20]~q ;
wire \regs[20][20]~q ;
wire \rfif.rdat1[20]~224_combout ;
wire \rfif.rdat1[20]~225_combout ;
wire \regs[18][20]~q ;
wire \regs[22][20]~q ;
wire \rfif.rdat1[20]~222_combout ;
wire \regs[26][20]~q ;
wire \regs[30][20]~q ;
wire \rfif.rdat1[20]~223_combout ;
wire \rfif.rdat1[20]~226_combout ;
wire \regs[10][20]~q ;
wire \regs[8][20]~q ;
wire \rfif.rdat1[20]~232_combout ;
wire \regs[9][20]~q ;
wire \rfif.rdat1[20]~233_combout ;
wire \regs[3][20]~q ;
wire \regs[1][20]~q ;
wire \regs[0][20]~q ;
wire \regs[2][20]~feeder_combout ;
wire \regs[2][20]~q ;
wire \rfif.rdat1[20]~234_combout ;
wire \rfif.rdat1[20]~235_combout ;
wire \rfif.rdat1[20]~236_combout ;
wire \regs[15][20]~q ;
wire \regs[13][20]~q ;
wire \rfif.rdat1[20]~237_combout ;
wire \regs[14][20]~feeder_combout ;
wire \regs[14][20]~q ;
wire \rfif.rdat1[20]~238_combout ;
wire \regs[6][20]~feeder_combout ;
wire \regs[6][20]~q ;
wire \regs[7][20]~q ;
wire \regs[5][20]~q ;
wire \rfif.rdat1[20]~230_combout ;
wire \rfif.rdat1[20]~231_combout ;
wire \rfif.rdat2[20]~238_combout ;
wire \rfif.rdat2[20]~239_combout ;
wire \rfif.rdat2[20]~233_combout ;
wire \rfif.rdat2[20]~234_combout ;
wire \regs[28][20]~q ;
wire \rfif.rdat2[20]~236_combout ;
wire \rfif.rdat2[20]~237_combout ;
wire \rfif.rdat2[20]~231_combout ;
wire \rfif.rdat2[20]~232_combout ;
wire \rfif.rdat2[20]~240_combout ;
wire \rfif.rdat2[20]~245_combout ;
wire \rfif.rdat2[20]~246_combout ;
wire \rfif.rdat2[20]~243_combout ;
wire \regs[11][20]~q ;
wire \rfif.rdat2[20]~244_combout ;
wire \rfif.rdat2[20]~247_combout ;
wire \regs[4][20]~q ;
wire \rfif.rdat2[20]~241_combout ;
wire \rfif.rdat2[20]~242_combout ;
wire \regs[12][20]~q ;
wire \rfif.rdat2[20]~248_combout ;
wire \rfif.rdat2[20]~249_combout ;
wire \rfif.rdat2[20]~250_combout ;
wire \regs[26][19]~q ;
wire \regs[18][19]~q ;
wire \rfif.rdat1[19]~240_combout ;
wire \regs[30][19]~q ;
wire \regs[22][19]~q ;
wire \rfif.rdat1[19]~241_combout ;
wire \regs[19][19]~q ;
wire \regs[23][19]~feeder_combout ;
wire \regs[23][19]~q ;
wire \rfif.rdat1[19]~247_combout ;
wire \regs[27][19]~q ;
wire \regs[31][19]~q ;
wire \rfif.rdat1[19]~248_combout ;
wire \regs[20][19]~q ;
wire \regs[28][19]~feeder_combout ;
wire \regs[28][19]~q ;
wire \rfif.rdat1[19]~245_combout ;
wire \regs[25][19]~q ;
wire \regs[29][19]~q ;
wire \rfif.rdat1[19]~243_combout ;
wire \rfif.rdat1[19]~246_combout ;
wire \regs[3][19]~feeder_combout ;
wire \regs[3][19]~q ;
wire \regs[0][19]~feeder_combout ;
wire \regs[0][19]~q ;
wire \rfif.rdat1[19]~254_combout ;
wire \rfif.rdat1[19]~255_combout ;
wire \regs[5][19]~feeder_combout ;
wire \regs[5][19]~q ;
wire \regs[7][19]~feeder_combout ;
wire \regs[7][19]~q ;
wire \rfif.rdat1[19]~253_combout ;
wire \rfif.rdat1[19]~256_combout ;
wire \regs[9][19]~feeder_combout ;
wire \regs[9][19]~q ;
wire \rfif.rdat1[19]~250_combout ;
wire \regs[11][19]~q ;
wire \regs[10][19]~q ;
wire \rfif.rdat1[19]~251_combout ;
wire \regs[15][19]~q ;
wire \regs[13][19]~feeder_combout ;
wire \regs[13][19]~q ;
wire \regs[14][19]~q ;
wire \regs[12][19]~q ;
wire \rfif.rdat1[19]~257_combout ;
wire \rfif.rdat1[19]~258_combout ;
wire \rfif.rdat2[19]~266_combout ;
wire \rfif.rdat2[19]~267_combout ;
wire \regs[4][19]~q ;
wire \regs[6][19]~q ;
wire \rfif.rdat2[19]~264_combout ;
wire \rfif.rdat2[19]~265_combout ;
wire \rfif.rdat2[19]~268_combout ;
wire \regs[8][19]~q ;
wire \rfif.rdat2[19]~262_combout ;
wire \rfif.rdat2[19]~263_combout ;
wire \rfif.rdat2[19]~270_combout ;
wire \rfif.rdat2[19]~271_combout ;
wire \rfif.rdat2[19]~252_combout ;
wire \rfif.rdat2[19]~253_combout ;
wire \rfif.rdat2[19]~259_combout ;
wire \rfif.rdat2[19]~260_combout ;
wire \regs[17][19]~q ;
wire \regs[21][19]~q ;
wire \rfif.rdat2[19]~254_combout ;
wire \rfif.rdat2[19]~255_combout ;
wire \regs[24][19]~q ;
wire \regs[16][19]~q ;
wire \rfif.rdat2[19]~256_combout ;
wire \rfif.rdat2[19]~257_combout ;
wire \rfif.rdat2[19]~258_combout ;
wire \rfif.rdat2[19]~261_combout ;
wire \regs[21][18]~q ;
wire \regs[29][18]~q ;
wire \regs[17][18]~q ;
wire \regs[25][18]~q ;
wire \rfif.rdat1[18]~260_combout ;
wire \rfif.rdat1[18]~261_combout ;
wire \regs[19][18]~feeder_combout ;
wire \regs[19][18]~q ;
wire \regs[27][18]~feeder_combout ;
wire \regs[27][18]~q ;
wire \rfif.rdat1[18]~267_combout ;
wire \regs[23][18]~q ;
wire \regs[31][18]~q ;
wire \rfif.rdat1[18]~268_combout ;
wire \regs[24][18]~q ;
wire \regs[20][18]~q ;
wire \rfif.rdat1[18]~264_combout ;
wire \rfif.rdat1[18]~265_combout ;
wire \regs[26][18]~q ;
wire \regs[22][18]~q ;
wire \rfif.rdat1[18]~262_combout ;
wire \rfif.rdat1[18]~263_combout ;
wire \rfif.rdat1[18]~266_combout ;
wire \regs[15][18]~q ;
wire \regs[14][18]~feeder_combout ;
wire \regs[14][18]~q ;
wire \regs[12][18]~q ;
wire \regs[13][18]~q ;
wire \rfif.rdat1[18]~277_combout ;
wire \rfif.rdat1[18]~278_combout ;
wire \regs[7][18]~q ;
wire \regs[6][18]~q ;
wire \regs[5][18]~q ;
wire \rfif.rdat1[18]~270_combout ;
wire \rfif.rdat1[18]~271_combout ;
wire \regs[11][18]~q ;
wire \regs[9][18]~q ;
wire \regs[10][18]~feeder_combout ;
wire \regs[10][18]~q ;
wire \rfif.rdat1[18]~272_combout ;
wire \rfif.rdat1[18]~273_combout ;
wire \regs[1][18]~feeder_combout ;
wire \regs[1][18]~q ;
wire \regs[3][18]~feeder_combout ;
wire \regs[3][18]~q ;
wire \regs[2][18]~q ;
wire \regs[0][18]~q ;
wire \rfif.rdat1[18]~274_combout ;
wire \rfif.rdat1[18]~275_combout ;
wire \rfif.rdat1[18]~276_combout ;
wire \rfif.rdat2[18]~274_combout ;
wire \rfif.rdat2[18]~280_combout ;
wire \rfif.rdat2[18]~281_combout ;
wire \regs[16][18]~q ;
wire \rfif.rdat2[18]~277_combout ;
wire \regs[28][18]~q ;
wire \rfif.rdat2[18]~278_combout ;
wire \regs[30][18]~q ;
wire \regs[18][18]~q ;
wire \rfif.rdat2[18]~275_combout ;
wire \rfif.rdat2[18]~276_combout ;
wire \rfif.rdat2[18]~279_combout ;
wire \rfif.rdat2[18]~282_combout ;
wire \regs[8][18]~q ;
wire \rfif.rdat2[18]~285_combout ;
wire \rfif.rdat2[18]~286_combout ;
wire \rfif.rdat2[18]~287_combout ;
wire \rfif.rdat2[18]~288_combout ;
wire \rfif.rdat2[18]~289_combout ;
wire \regs[4][18]~q ;
wire \rfif.rdat2[18]~283_combout ;
wire \rfif.rdat2[18]~284_combout ;
wire \rfif.rdat2[18]~290_combout ;
wire \rfif.rdat2[18]~291_combout ;
wire \rfif.rdat2[18]~292_combout ;
wire \regs[18][17]~q ;
wire \regs[26][17]~q ;
wire \rfif.rdat1[17]~280_combout ;
wire \regs[30][17]~q ;
wire \regs[22][17]~q ;
wire \rfif.rdat1[17]~281_combout ;
wire \regs[21][17]~q ;
wire \rfif.rdat1[17]~282_combout ;
wire \regs[25][17]~q ;
wire \regs[29][17]~q ;
wire \rfif.rdat1[17]~283_combout ;
wire \regs[20][17]~q ;
wire \regs[28][17]~q ;
wire \rfif.rdat1[17]~285_combout ;
wire \rfif.rdat1[17]~286_combout ;
wire \regs[27][17]~feeder_combout ;
wire \regs[27][17]~q ;
wire \regs[23][17]~q ;
wire \regs[19][17]~q ;
wire \rfif.rdat1[17]~287_combout ;
wire \regs[31][17]~feeder_combout ;
wire \regs[31][17]~q ;
wire \rfif.rdat1[17]~288_combout ;
wire \regs[13][17]~q ;
wire \regs[15][17]~feeder_combout ;
wire \regs[15][17]~q ;
wire \regs[12][17]~q ;
wire \rfif.rdat1[17]~297_combout ;
wire \rfif.rdat1[17]~298_combout ;
wire \regs[9][17]~q ;
wire \regs[8][17]~q ;
wire \rfif.rdat1[17]~290_combout ;
wire \regs[11][17]~q ;
wire \regs[10][17]~q ;
wire \rfif.rdat1[17]~291_combout ;
wire \regs[1][17]~q ;
wire \regs[0][17]~q ;
wire \rfif.rdat1[17]~294_combout ;
wire \regs[3][17]~feeder_combout ;
wire \regs[3][17]~q ;
wire \rfif.rdat1[17]~295_combout ;
wire \regs[7][17]~q ;
wire \regs[5][17]~q ;
wire \rfif.rdat1[17]~293_combout ;
wire \rfif.rdat1[17]~296_combout ;
wire \regs[17][17]~q ;
wire \rfif.rdat2[17]~296_combout ;
wire \rfif.rdat2[17]~297_combout ;
wire \regs[24][17]~feeder_combout ;
wire \regs[24][17]~q ;
wire \rfif.rdat2[17]~298_combout ;
wire \rfif.rdat2[17]~299_combout ;
wire \rfif.rdat2[17]~300_combout ;
wire \rfif.rdat2[17]~301_combout ;
wire \rfif.rdat2[17]~302_combout ;
wire \rfif.rdat2[17]~294_combout ;
wire \rfif.rdat2[17]~295_combout ;
wire \rfif.rdat2[17]~303_combout ;
wire \rfif.rdat2[17]~304_combout ;
wire \rfif.rdat2[17]~305_combout ;
wire \regs[14][17]~feeder_combout ;
wire \regs[14][17]~q ;
wire \rfif.rdat2[17]~311_combout ;
wire \rfif.rdat2[17]~312_combout ;
wire \regs[4][17]~q ;
wire \regs[6][17]~feeder_combout ;
wire \regs[6][17]~q ;
wire \rfif.rdat2[17]~306_combout ;
wire \rfif.rdat2[17]~307_combout ;
wire \rfif.rdat2[17]~310_combout ;
wire \rfif.rdat2[17]~313_combout ;
wire \regs[31][16]~q ;
wire \regs[23][16]~q ;
wire \regs[27][16]~feeder_combout ;
wire \regs[27][16]~q ;
wire \regs[19][16]~feeder_combout ;
wire \regs[19][16]~q ;
wire \rfif.rdat1[16]~307_combout ;
wire \rfif.rdat1[16]~308_combout ;
wire \regs[24][16]~q ;
wire \regs[28][16]~q ;
wire \rfif.rdat1[16]~305_combout ;
wire \regs[26][16]~q ;
wire \regs[30][16]~q ;
wire \rfif.rdat1[16]~303_combout ;
wire \rfif.rdat1[16]~306_combout ;
wire \regs[25][16]~q ;
wire \regs[17][16]~q ;
wire \rfif.rdat1[16]~300_combout ;
wire \regs[29][16]~q ;
wire \regs[21][16]~q ;
wire \rfif.rdat1[16]~301_combout ;
wire \regs[10][16]~q ;
wire \regs[8][16]~q ;
wire \rfif.rdat1[16]~312_combout ;
wire \regs[9][16]~q ;
wire \rfif.rdat1[16]~313_combout ;
wire \regs[1][16]~feeder_combout ;
wire \regs[1][16]~q ;
wire \regs[2][16]~q ;
wire \rfif.rdat1[16]~314_combout ;
wire \rfif.rdat1[16]~315_combout ;
wire \rfif.rdat1[16]~316_combout ;
wire \regs[7][16]~q ;
wire \regs[6][16]~q ;
wire \regs[5][16]~q ;
wire \rfif.rdat1[16]~310_combout ;
wire \rfif.rdat1[16]~311_combout ;
wire \regs[15][16]~feeder_combout ;
wire \regs[15][16]~q ;
wire \regs[13][16]~q ;
wire \rfif.rdat1[16]~317_combout ;
wire \regs[14][16]~feeder_combout ;
wire \regs[14][16]~q ;
wire \rfif.rdat1[16]~318_combout ;
wire \regs[12][16]~q ;
wire \rfif.rdat2[16]~332_combout ;
wire \rfif.rdat2[16]~333_combout ;
wire \regs[0][16]~q ;
wire \rfif.rdat2[16]~329_combout ;
wire \rfif.rdat2[16]~330_combout ;
wire \regs[11][16]~q ;
wire \rfif.rdat2[16]~328_combout ;
wire \rfif.rdat2[16]~331_combout ;
wire \regs[4][16]~q ;
wire \rfif.rdat2[16]~325_combout ;
wire \rfif.rdat2[16]~326_combout ;
wire \rfif.rdat2[16]~334_combout ;
wire \rfif.rdat2[16]~322_combout ;
wire \rfif.rdat2[16]~323_combout ;
wire \rfif.rdat2[16]~320_combout ;
wire \rfif.rdat2[16]~321_combout ;
wire \rfif.rdat2[16]~315_combout ;
wire \rfif.rdat2[16]~316_combout ;
wire \rfif.rdat2[16]~324_combout ;
wire \regs[26][15]~q ;
wire \rfif.rdat1[15]~320_combout ;
wire \regs[30][15]~q ;
wire \regs[22][15]~q ;
wire \rfif.rdat1[15]~321_combout ;
wire \regs[20][15]~q ;
wire \regs[24][15]~q ;
wire \regs[16][15]~q ;
wire \rfif.rdat1[15]~324_combout ;
wire \rfif.rdat1[15]~325_combout ;
wire \regs[21][15]~q ;
wire \regs[17][15]~q ;
wire \rfif.rdat1[15]~322_combout ;
wire \regs[25][15]~q ;
wire \regs[29][15]~q ;
wire \rfif.rdat1[15]~323_combout ;
wire \rfif.rdat1[15]~326_combout ;
wire \regs[31][15]~q ;
wire \regs[27][15]~feeder_combout ;
wire \regs[27][15]~q ;
wire \regs[23][15]~q ;
wire \regs[19][15]~q ;
wire \rfif.rdat1[15]~327_combout ;
wire \rfif.rdat1[15]~328_combout ;
wire \regs[10][15]~q ;
wire \regs[11][15]~q ;
wire \regs[9][15]~q ;
wire \regs[8][15]~q ;
wire \rfif.rdat1[15]~330_combout ;
wire \rfif.rdat1[15]~331_combout ;
wire \regs[7][15]~q ;
wire \regs[5][15]~q ;
wire \rfif.rdat1[15]~333_combout ;
wire \regs[2][15]~q ;
wire \regs[3][15]~q ;
wire \regs[1][15]~q ;
wire \regs[0][15]~q ;
wire \rfif.rdat1[15]~334_combout ;
wire \rfif.rdat1[15]~335_combout ;
wire \rfif.rdat1[15]~336_combout ;
wire \regs[12][15]~q ;
wire \regs[14][15]~q ;
wire \rfif.rdat1[15]~337_combout ;
wire \regs[13][15]~q ;
wire \regs[15][15]~feeder_combout ;
wire \regs[15][15]~q ;
wire \rfif.rdat1[15]~338_combout ;
wire \rfif.rdat2[15]~346_combout ;
wire \rfif.rdat2[15]~347_combout ;
wire \rfif.rdat2[15]~353_combout ;
wire \rfif.rdat2[15]~354_combout ;
wire \rfif.rdat2[15]~350_combout ;
wire \rfif.rdat2[15]~351_combout ;
wire \regs[4][15]~q ;
wire \regs[6][15]~q ;
wire \rfif.rdat2[15]~348_combout ;
wire \rfif.rdat2[15]~349_combout ;
wire \rfif.rdat2[15]~352_combout ;
wire \rfif.rdat2[15]~355_combout ;
wire \rfif.rdat2[15]~344_combout ;
wire \regs[18][15]~q ;
wire \rfif.rdat2[15]~336_combout ;
wire \rfif.rdat2[15]~337_combout ;
wire \rfif.rdat2[15]~338_combout ;
wire \rfif.rdat2[15]~339_combout ;
wire \regs[28][15]~q ;
wire \rfif.rdat2[15]~340_combout ;
wire \rfif.rdat2[15]~341_combout ;
wire \rfif.rdat2[15]~342_combout ;
wire \rfif.rdat2[15]~345_combout ;
wire \regs[17][14]~q ;
wire \regs[25][14]~q ;
wire \rfif.rdat1[14]~340_combout ;
wire \regs[29][14]~q ;
wire \regs[21][14]~q ;
wire \rfif.rdat1[14]~341_combout ;
wire \regs[31][14]~q ;
wire \regs[23][14]~q ;
wire \regs[27][14]~q ;
wire \regs[19][14]~q ;
wire \rfif.rdat1[14]~347_combout ;
wire \rfif.rdat1[14]~348_combout ;
wire \regs[24][14]~q ;
wire \regs[28][14]~q ;
wire \rfif.rdat1[14]~345_combout ;
wire \regs[30][14]~q ;
wire \regs[26][14]~q ;
wire \regs[18][14]~q ;
wire \regs[22][14]~q ;
wire \rfif.rdat1[14]~342_combout ;
wire \rfif.rdat1[14]~343_combout ;
wire \rfif.rdat1[14]~346_combout ;
wire \regs[13][14]~q ;
wire \rfif.rdat1[14]~357_combout ;
wire \regs[14][14]~q ;
wire \regs[15][14]~q ;
wire \rfif.rdat1[14]~358_combout ;
wire \regs[7][14]~q ;
wire \regs[6][14]~q ;
wire \regs[4][14]~q ;
wire \rfif.rdat1[14]~350_combout ;
wire \rfif.rdat1[14]~351_combout ;
wire \regs[11][14]~feeder_combout ;
wire \regs[11][14]~q ;
wire \regs[9][14]~feeder_combout ;
wire \regs[9][14]~q ;
wire \regs[8][14]~q ;
wire \regs[10][14]~q ;
wire \rfif.rdat1[14]~352_combout ;
wire \rfif.rdat1[14]~353_combout ;
wire \regs[1][14]~q ;
wire \regs[2][14]~q ;
wire \rfif.rdat1[14]~354_combout ;
wire \rfif.rdat1[14]~355_combout ;
wire \rfif.rdat1[14]~356_combout ;
wire \rfif.rdat2[14]~358_combout ;
wire \regs[20][14]~q ;
wire \rfif.rdat2[14]~361_combout ;
wire \rfif.rdat2[14]~362_combout ;
wire \rfif.rdat2[14]~359_combout ;
wire \rfif.rdat2[14]~360_combout ;
wire \rfif.rdat2[14]~363_combout ;
wire \rfif.rdat2[14]~364_combout ;
wire \rfif.rdat2[14]~365_combout ;
wire \rfif.rdat2[14]~366_combout ;
wire \regs[5][14]~q ;
wire \rfif.rdat2[14]~367_combout ;
wire \rfif.rdat2[14]~368_combout ;
wire \regs[12][14]~q ;
wire \rfif.rdat2[14]~374_combout ;
wire \rfif.rdat2[14]~375_combout ;
wire \rfif.rdat2[14]~369_combout ;
wire \rfif.rdat2[14]~370_combout ;
wire \regs[0][14]~q ;
wire \rfif.rdat2[14]~371_combout ;
wire \regs[3][14]~feeder_combout ;
wire \regs[3][14]~q ;
wire \rfif.rdat2[14]~372_combout ;
wire \rfif.rdat2[14]~373_combout ;
wire \rfif.rdat2[14]~376_combout ;
wire \regs[18][13]~q ;
wire \regs[26][13]~q ;
wire \rfif.rdat2[13]~378_combout ;
wire \regs[22][13]~q ;
wire \regs[30][13]~q ;
wire \rfif.rdat2[13]~379_combout ;
wire \regs[25][13]~q ;
wire \regs[29][13]~q ;
wire \regs[17][13]~q ;
wire \regs[21][13]~feeder_combout ;
wire \regs[21][13]~q ;
wire \rfif.rdat2[13]~380_combout ;
wire \rfif.rdat2[13]~381_combout ;
wire \rfif.rdat2[13]~384_combout ;
wire \regs[27][13]~feeder_combout ;
wire \regs[27][13]~q ;
wire \regs[23][13]~feeder_combout ;
wire \regs[23][13]~q ;
wire \regs[19][13]~q ;
wire \rfif.rdat2[13]~385_combout ;
wire \rfif.rdat2[13]~386_combout ;
wire \rfif.rdat2[13]~387_combout ;
wire \regs[2][13]~q ;
wire \regs[0][13]~q ;
wire \regs[1][13]~feeder_combout ;
wire \regs[1][13]~q ;
wire \rfif.rdat2[13]~392_combout ;
wire \rfif.rdat2[13]~393_combout ;
wire \rfif.rdat2[13]~394_combout ;
wire \regs[13][13]~q ;
wire \regs[15][13]~feeder_combout ;
wire \regs[15][13]~q ;
wire \regs[12][13]~q ;
wire \regs[14][13]~feeder_combout ;
wire \regs[14][13]~q ;
wire \rfif.rdat2[13]~395_combout ;
wire \rfif.rdat2[13]~396_combout ;
wire \regs[10][13]~q ;
wire \regs[11][13]~feeder_combout ;
wire \regs[11][13]~q ;
wire \regs[8][13]~q ;
wire \regs[9][13]~feeder_combout ;
wire \regs[9][13]~q ;
wire \rfif.rdat2[13]~388_combout ;
wire \rfif.rdat2[13]~389_combout ;
wire \rfif.rdat2[13]~397_combout ;
wire \rfif.rdat1[13]~362_combout ;
wire \rfif.rdat1[13]~363_combout ;
wire \regs[28][13]~q ;
wire \regs[24][13]~q ;
wire \rfif.rdat1[13]~365_combout ;
wire \rfif.rdat1[13]~366_combout ;
wire \rfif.rdat1[13]~360_combout ;
wire \rfif.rdat1[13]~361_combout ;
wire \rfif.rdat1[13]~367_combout ;
wire \regs[31][13]~feeder_combout ;
wire \regs[31][13]~q ;
wire \rfif.rdat1[13]~368_combout ;
wire \regs[7][13]~feeder_combout ;
wire \regs[7][13]~q ;
wire \regs[6][13]~q ;
wire \regs[5][13]~q ;
wire \rfif.rdat1[13]~370_combout ;
wire \rfif.rdat1[13]~371_combout ;
wire \rfif.rdat1[13]~377_combout ;
wire \rfif.rdat1[13]~378_combout ;
wire \rfif.rdat1[13]~374_combout ;
wire \regs[3][13]~feeder_combout ;
wire \regs[3][13]~q ;
wire \rfif.rdat1[13]~375_combout ;
wire \rfif.rdat1[13]~372_combout ;
wire \rfif.rdat1[13]~373_combout ;
wire \rfif.rdat1[13]~376_combout ;
wire \regs[21][12]~q ;
wire \regs[25][12]~q ;
wire \rfif.rdat2[12]~399_combout ;
wire \rfif.rdat2[12]~400_combout ;
wire \regs[28][12]~q ;
wire \regs[16][12]~q ;
wire \regs[20][12]~q ;
wire \rfif.rdat2[12]~403_combout ;
wire \rfif.rdat2[12]~404_combout ;
wire \regs[26][12]~q ;
wire \regs[30][12]~q ;
wire \regs[18][12]~q ;
wire \regs[22][12]~q ;
wire \rfif.rdat2[12]~401_combout ;
wire \rfif.rdat2[12]~402_combout ;
wire \rfif.rdat2[12]~405_combout ;
wire \regs[23][12]~q ;
wire \regs[31][12]~q ;
wire \rfif.rdat2[12]~407_combout ;
wire \rfif.rdat2[12]~408_combout ;
wire \regs[6][12]~q ;
wire \regs[4][12]~q ;
wire \rfif.rdat2[12]~409_combout ;
wire \rfif.rdat2[12]~410_combout ;
wire \regs[0][12]~q ;
wire \rfif.rdat2[12]~413_combout ;
wire \regs[3][12]~q ;
wire \regs[1][12]~q ;
wire \rfif.rdat2[12]~414_combout ;
wire \regs[8][12]~q ;
wire \regs[10][12]~feeder_combout ;
wire \regs[10][12]~q ;
wire \rfif.rdat2[12]~411_combout ;
wire \regs[11][12]~q ;
wire \regs[9][12]~q ;
wire \rfif.rdat2[12]~412_combout ;
wire \rfif.rdat2[12]~415_combout ;
wire \regs[15][12]~feeder_combout ;
wire \regs[15][12]~q ;
wire \regs[14][12]~feeder_combout ;
wire \regs[14][12]~q ;
wire \rfif.rdat2[12]~417_combout ;
wire \rfif.rdat2[12]~418_combout ;
wire \regs[24][12]~q ;
wire \rfif.rdat1[12]~384_combout ;
wire \rfif.rdat1[12]~385_combout ;
wire \regs[29][12]~q ;
wire \regs[17][12]~q ;
wire \rfif.rdat1[12]~382_combout ;
wire \rfif.rdat1[12]~383_combout ;
wire \rfif.rdat1[12]~386_combout ;
wire \rfif.rdat1[12]~387_combout ;
wire \regs[27][12]~q ;
wire \rfif.rdat1[12]~388_combout ;
wire \rfif.rdat1[12]~380_combout ;
wire \rfif.rdat1[12]~381_combout ;
wire \rfif.rdat1[12]~390_combout ;
wire \rfif.rdat1[12]~391_combout ;
wire \regs[2][12]~q ;
wire \rfif.rdat1[12]~395_combout ;
wire \regs[5][12]~feeder_combout ;
wire \regs[5][12]~q ;
wire \rfif.rdat1[12]~392_combout ;
wire \rfif.rdat1[12]~393_combout ;
wire \rfif.rdat1[12]~396_combout ;
wire \regs[12][12]~q ;
wire \rfif.rdat1[12]~397_combout ;
wire \regs[13][12]~q ;
wire \rfif.rdat1[12]~398_combout ;
wire \regs[11][11]~feeder_combout ;
wire \regs[11][11]~q ;
wire \regs[10][11]~q ;
wire \regs[8][11]~q ;
wire \regs[9][11]~feeder_combout ;
wire \regs[9][11]~q ;
wire \rfif.rdat2[11]~430_combout ;
wire \rfif.rdat2[11]~431_combout ;
wire \regs[13][11]~q ;
wire \regs[12][11]~q ;
wire \regs[14][11]~q ;
wire \rfif.rdat2[11]~437_combout ;
wire \rfif.rdat2[11]~438_combout ;
wire \regs[4][11]~q ;
wire \rfif.rdat2[11]~432_combout ;
wire \regs[7][11]~q ;
wire \regs[5][11]~q ;
wire \rfif.rdat2[11]~433_combout ;
wire \rfif.rdat2[11]~436_combout ;
wire \rfif.rdat2[11]~439_combout ;
wire \regs[22][11]~q ;
wire \regs[18][11]~q ;
wire \regs[26][11]~q ;
wire \rfif.rdat2[11]~420_combout ;
wire \rfif.rdat2[11]~421_combout ;
wire \regs[27][11]~q ;
wire \regs[31][11]~q ;
wire \regs[19][11]~q ;
wire \regs[23][11]~q ;
wire \rfif.rdat2[11]~427_combout ;
wire \rfif.rdat2[11]~428_combout ;
wire \regs[28][11]~q ;
wire \regs[20][11]~q ;
wire \rfif.rdat2[11]~425_combout ;
wire \regs[25][11]~q ;
wire \regs[29][11]~q ;
wire \regs[17][11]~q ;
wire \regs[21][11]~q ;
wire \rfif.rdat2[11]~422_combout ;
wire \rfif.rdat2[11]~423_combout ;
wire \rfif.rdat2[11]~426_combout ;
wire \rfif.rdat2[11]~429_combout ;
wire \rfif.rdat1[11]~407_combout ;
wire \rfif.rdat1[11]~408_combout ;
wire \rfif.rdat1[11]~400_combout ;
wire \rfif.rdat1[11]~401_combout ;
wire \rfif.rdat1[11]~404_combout ;
wire \regs[24][11]~q ;
wire \rfif.rdat1[11]~405_combout ;
wire \rfif.rdat1[11]~402_combout ;
wire \regs[30][11]~q ;
wire \rfif.rdat1[11]~403_combout ;
wire \rfif.rdat1[11]~406_combout ;
wire \rfif.rdat1[11]~417_combout ;
wire \regs[15][11]~q ;
wire \rfif.rdat1[11]~418_combout ;
wire \rfif.rdat1[11]~412_combout ;
wire \rfif.rdat1[11]~413_combout ;
wire \regs[2][11]~q ;
wire \regs[0][11]~q ;
wire \rfif.rdat1[11]~414_combout ;
wire \regs[1][11]~q ;
wire \regs[3][11]~q ;
wire \rfif.rdat1[11]~415_combout ;
wire \rfif.rdat1[11]~416_combout ;
wire \regs[6][11]~q ;
wire \rfif.rdat1[11]~410_combout ;
wire \rfif.rdat1[11]~411_combout ;
wire \regs[13][10]~q ;
wire \regs[12][10]~q ;
wire \rfif.rdat2[10]~458_combout ;
wire \regs[14][10]~q ;
wire \regs[15][10]~feeder_combout ;
wire \regs[15][10]~q ;
wire \rfif.rdat2[10]~459_combout ;
wire \regs[6][10]~q ;
wire \regs[7][10]~q ;
wire \regs[4][10]~q ;
wire \regs[5][10]~q ;
wire \rfif.rdat2[10]~451_combout ;
wire \rfif.rdat2[10]~452_combout ;
wire \regs[9][10]~q ;
wire \regs[11][10]~q ;
wire \regs[8][10]~q ;
wire \regs[10][10]~q ;
wire \rfif.rdat2[10]~453_combout ;
wire \rfif.rdat2[10]~454_combout ;
wire \rfif.rdat2[10]~457_combout ;
wire \rfif.rdat2[10]~460_combout ;
wire \regs[25][10]~q ;
wire \regs[17][10]~q ;
wire \rfif.rdat2[10]~441_combout ;
wire \regs[21][10]~q ;
wire \regs[29][10]~q ;
wire \rfif.rdat2[10]~442_combout ;
wire \regs[19][10]~q ;
wire \regs[27][10]~feeder_combout ;
wire \regs[27][10]~q ;
wire \rfif.rdat2[10]~448_combout ;
wire \regs[23][10]~q ;
wire \rfif.rdat2[10]~449_combout ;
wire \regs[28][10]~q ;
wire \regs[16][10]~q ;
wire \regs[20][10]~q ;
wire \rfif.rdat2[10]~445_combout ;
wire \rfif.rdat2[10]~446_combout ;
wire \regs[18][10]~q ;
wire \regs[22][10]~q ;
wire \rfif.rdat2[10]~443_combout ;
wire \regs[30][10]~q ;
wire \regs[26][10]~q ;
wire \rfif.rdat2[10]~444_combout ;
wire \rfif.rdat2[10]~447_combout ;
wire \rfif.rdat2[10]~450_combout ;
wire \rfif.rdat1[10]~427_combout ;
wire \regs[31][10]~feeder_combout ;
wire \regs[31][10]~q ;
wire \rfif.rdat1[10]~428_combout ;
wire \rfif.rdat1[10]~420_combout ;
wire \rfif.rdat1[10]~421_combout ;
wire \regs[24][10]~q ;
wire \rfif.rdat1[10]~424_combout ;
wire \rfif.rdat1[10]~425_combout ;
wire \rfif.rdat1[10]~422_combout ;
wire \rfif.rdat1[10]~423_combout ;
wire \rfif.rdat1[10]~426_combout ;
wire \rfif.rdat1[10]~437_combout ;
wire \rfif.rdat1[10]~438_combout ;
wire \rfif.rdat1[10]~433_combout ;
wire \regs[3][10]~q ;
wire \regs[2][10]~q ;
wire \rfif.rdat1[10]~435_combout ;
wire \rfif.rdat1[10]~436_combout ;
wire \rfif.rdat1[10]~430_combout ;
wire \rfif.rdat1[10]~431_combout ;
wire \regs[25][9]~q ;
wire \regs[29][9]~q ;
wire \rfif.rdat2[9]~465_combout ;
wire \regs[28][9]~q ;
wire \regs[16][9]~q ;
wire \regs[24][9]~q ;
wire \rfif.rdat2[9]~466_combout ;
wire \rfif.rdat2[9]~467_combout ;
wire \rfif.rdat2[9]~468_combout ;
wire \regs[22][9]~q ;
wire \regs[30][9]~q ;
wire \rfif.rdat2[9]~463_combout ;
wire \regs[31][9]~q ;
wire \regs[23][9]~q ;
wire \regs[19][9]~q ;
wire \rfif.rdat2[9]~469_combout ;
wire \rfif.rdat2[9]~470_combout ;
wire \rfif.rdat2[9]~471_combout ;
wire \regs[11][9]~feeder_combout ;
wire \regs[11][9]~q ;
wire \regs[10][9]~q ;
wire \rfif.rdat2[9]~473_combout ;
wire \regs[13][9]~q ;
wire \regs[12][9]~q ;
wire \regs[14][9]~q ;
wire \rfif.rdat2[9]~479_combout ;
wire \rfif.rdat2[9]~480_combout ;
wire \regs[2][9]~q ;
wire \regs[3][9]~q ;
wire \regs[0][9]~q ;
wire \rfif.rdat2[9]~476_combout ;
wire \rfif.rdat2[9]~477_combout ;
wire \regs[5][9]~q ;
wire \regs[7][9]~q ;
wire \regs[4][9]~q ;
wire \regs[6][9]~q ;
wire \rfif.rdat2[9]~474_combout ;
wire \rfif.rdat2[9]~475_combout ;
wire \rfif.rdat2[9]~478_combout ;
wire \rfif.rdat2[9]~481_combout ;
wire \regs[21][9]~q ;
wire \regs[17][9]~q ;
wire \rfif.rdat1[9]~440_combout ;
wire \rfif.rdat1[9]~441_combout ;
wire \regs[27][9]~q ;
wire \rfif.rdat1[9]~447_combout ;
wire \rfif.rdat1[9]~448_combout ;
wire \rfif.rdat1[9]~445_combout ;
wire \regs[26][9]~q ;
wire \regs[18][9]~q ;
wire \rfif.rdat1[9]~442_combout ;
wire \rfif.rdat1[9]~443_combout ;
wire \rfif.rdat1[9]~446_combout ;
wire \regs[1][9]~q ;
wire \rfif.rdat1[9]~455_combout ;
wire \rfif.rdat1[9]~452_combout ;
wire \rfif.rdat1[9]~453_combout ;
wire \rfif.rdat1[9]~456_combout ;
wire \regs[15][9]~q ;
wire \rfif.rdat1[9]~457_combout ;
wire \rfif.rdat1[9]~458_combout ;
wire \rfif.rdat1[9]~450_combout ;
wire \rfif.rdat1[9]~451_combout ;
wire \regs[25][8]~q ;
wire \regs[17][8]~q ;
wire \rfif.rdat2[8]~483_combout ;
wire \regs[21][8]~q ;
wire \regs[29][8]~q ;
wire \rfif.rdat2[8]~484_combout ;
wire \regs[31][8]~feeder_combout ;
wire \regs[31][8]~q ;
wire \regs[19][8]~q ;
wire \regs[27][8]~feeder_combout ;
wire \regs[27][8]~q ;
wire \rfif.rdat2[8]~490_combout ;
wire \rfif.rdat2[8]~491_combout ;
wire \regs[30][8]~q ;
wire \regs[26][8]~q ;
wire \rfif.rdat2[8]~486_combout ;
wire \rfif.rdat2[8]~489_combout ;
wire \rfif.rdat2[8]~492_combout ;
wire \regs[7][8]~feeder_combout ;
wire \regs[7][8]~q ;
wire \regs[4][8]~q ;
wire \regs[5][8]~feeder_combout ;
wire \regs[5][8]~q ;
wire \rfif.rdat2[8]~493_combout ;
wire \regs[6][8]~feeder_combout ;
wire \regs[6][8]~q ;
wire \rfif.rdat2[8]~494_combout ;
wire \regs[15][8]~feeder_combout ;
wire \regs[15][8]~q ;
wire \regs[12][8]~q ;
wire \regs[13][8]~q ;
wire \rfif.rdat2[8]~500_combout ;
wire \regs[14][8]~feeder_combout ;
wire \regs[14][8]~q ;
wire \rfif.rdat2[8]~501_combout ;
wire \regs[1][8]~q ;
wire \regs[3][8]~q ;
wire \regs[0][8]~q ;
wire \regs[2][8]~feeder_combout ;
wire \regs[2][8]~q ;
wire \rfif.rdat2[8]~497_combout ;
wire \rfif.rdat2[8]~498_combout ;
wire \regs[9][8]~q ;
wire \regs[11][8]~q ;
wire \regs[10][8]~q ;
wire \regs[8][8]~feeder_combout ;
wire \regs[8][8]~q ;
wire \rfif.rdat2[8]~495_combout ;
wire \rfif.rdat2[8]~496_combout ;
wire \rfif.rdat2[8]~499_combout ;
wire \rfif.rdat2[8]~502_combout ;
wire \regs[18][8]~q ;
wire \rfif.rdat1[8]~460_combout ;
wire \regs[22][8]~q ;
wire \rfif.rdat1[8]~461_combout ;
wire \rfif.rdat1[8]~462_combout ;
wire \rfif.rdat1[8]~463_combout ;
wire \regs[28][8]~feeder_combout ;
wire \regs[28][8]~q ;
wire \regs[20][8]~feeder_combout ;
wire \regs[20][8]~q ;
wire \rfif.rdat1[8]~465_combout ;
wire \rfif.rdat1[8]~466_combout ;
wire \regs[23][8]~q ;
wire \rfif.rdat1[8]~467_combout ;
wire \rfif.rdat1[8]~468_combout ;
wire \rfif.rdat1[8]~470_combout ;
wire \rfif.rdat1[8]~471_combout ;
wire \rfif.rdat1[8]~477_combout ;
wire \rfif.rdat1[8]~478_combout ;
wire \rfif.rdat1[8]~472_combout ;
wire \rfif.rdat1[8]~473_combout ;
wire \rfif.rdat1[8]~474_combout ;
wire \rfif.rdat1[8]~475_combout ;
wire \rfif.rdat1[8]~476_combout ;
wire \regs[8][7]~q ;
wire \regs[9][7]~feeder_combout ;
wire \regs[9][7]~q ;
wire \rfif.rdat2[7]~514_combout ;
wire \regs[11][7]~q ;
wire \rfif.rdat2[7]~515_combout ;
wire \regs[12][7]~q ;
wire \regs[14][7]~q ;
wire \rfif.rdat2[7]~521_combout ;
wire \regs[13][7]~feeder_combout ;
wire \regs[13][7]~q ;
wire \regs[15][7]~q ;
wire \rfif.rdat2[7]~522_combout ;
wire \regs[4][7]~q ;
wire \regs[6][7]~q ;
wire \rfif.rdat2[7]~516_combout ;
wire \regs[7][7]~q ;
wire \regs[5][7]~q ;
wire \rfif.rdat2[7]~517_combout ;
wire \regs[3][7]~feeder_combout ;
wire \regs[3][7]~q ;
wire \regs[2][7]~q ;
wire \regs[0][7]~q ;
wire \regs[1][7]~q ;
wire \rfif.rdat2[7]~518_combout ;
wire \rfif.rdat2[7]~519_combout ;
wire \rfif.rdat2[7]~520_combout ;
wire \rfif.rdat2[7]~523_combout ;
wire \regs[22][7]~q ;
wire \regs[18][7]~q ;
wire \regs[26][7]~q ;
wire \rfif.rdat2[7]~504_combout ;
wire \rfif.rdat2[7]~505_combout ;
wire \regs[19][7]~q ;
wire \regs[23][7]~q ;
wire \rfif.rdat2[7]~511_combout ;
wire \regs[31][7]~q ;
wire \regs[27][7]~q ;
wire \rfif.rdat2[7]~512_combout ;
wire \regs[25][7]~q ;
wire \regs[29][7]~q ;
wire \regs[17][7]~q ;
wire \regs[21][7]~q ;
wire \rfif.rdat2[7]~506_combout ;
wire \rfif.rdat2[7]~507_combout ;
wire \rfif.rdat2[7]~510_combout ;
wire \rfif.rdat2[7]~513_combout ;
wire \rfif.rdat1[7]~480_combout ;
wire \rfif.rdat1[7]~481_combout ;
wire \rfif.rdat1[7]~487_combout ;
wire \rfif.rdat1[7]~488_combout ;
wire \regs[20][7]~q ;
wire \rfif.rdat1[7]~484_combout ;
wire \regs[24][7]~q ;
wire \rfif.rdat1[7]~485_combout ;
wire \rfif.rdat1[7]~482_combout ;
wire \regs[30][7]~q ;
wire \rfif.rdat1[7]~483_combout ;
wire \rfif.rdat1[7]~486_combout ;
wire \regs[10][7]~q ;
wire \rfif.rdat1[7]~492_combout ;
wire \rfif.rdat1[7]~493_combout ;
wire \rfif.rdat1[7]~494_combout ;
wire \rfif.rdat1[7]~495_combout ;
wire \rfif.rdat1[7]~496_combout ;
wire \rfif.rdat1[7]~490_combout ;
wire \rfif.rdat1[7]~491_combout ;
wire \rfif.rdat1[7]~497_combout ;
wire \rfif.rdat1[7]~498_combout ;
wire \regs[26][6]~q ;
wire \regs[30][6]~q ;
wire \regs[22][6]~q ;
wire \regs[18][6]~q ;
wire \rfif.rdat2[6]~527_combout ;
wire \rfif.rdat2[6]~528_combout ;
wire \rfif.rdat2[6]~531_combout ;
wire \regs[21][6]~q ;
wire \regs[17][6]~q ;
wire \regs[25][6]~q ;
wire \rfif.rdat2[6]~525_combout ;
wire \rfif.rdat2[6]~526_combout ;
wire \regs[23][6]~q ;
wire \regs[31][6]~feeder_combout ;
wire \regs[31][6]~q ;
wire \rfif.rdat2[6]~533_combout ;
wire \rfif.rdat2[6]~534_combout ;
wire \regs[6][6]~q ;
wire \regs[5][6]~q ;
wire \regs[4][6]~q ;
wire \rfif.rdat2[6]~535_combout ;
wire \rfif.rdat2[6]~536_combout ;
wire \regs[15][6]~feeder_combout ;
wire \regs[15][6]~q ;
wire \regs[14][6]~q ;
wire \rfif.rdat2[6]~543_combout ;
wire \regs[1][6]~q ;
wire \regs[3][6]~q ;
wire \regs[0][6]~q ;
wire \rfif.rdat2[6]~539_combout ;
wire \rfif.rdat2[6]~540_combout ;
wire \regs[10][6]~q ;
wire \regs[8][6]~feeder_combout ;
wire \regs[8][6]~q ;
wire \rfif.rdat2[6]~537_combout ;
wire \regs[11][6]~q ;
wire \regs[9][6]~feeder_combout ;
wire \regs[9][6]~q ;
wire \rfif.rdat2[6]~538_combout ;
wire \rfif.rdat2[6]~541_combout ;
wire \rfif.rdat2[6]~544_combout ;
wire \rfif.rdat1[6]~500_combout ;
wire \rfif.rdat1[6]~501_combout ;
wire \regs[27][6]~feeder_combout ;
wire \regs[27][6]~q ;
wire \regs[19][6]~q ;
wire \rfif.rdat1[6]~507_combout ;
wire \rfif.rdat1[6]~508_combout ;
wire \regs[20][6]~feeder_combout ;
wire \regs[20][6]~q ;
wire \regs[28][6]~feeder_combout ;
wire \regs[28][6]~q ;
wire \rfif.rdat1[6]~505_combout ;
wire \rfif.rdat1[6]~502_combout ;
wire \regs[29][6]~q ;
wire \rfif.rdat1[6]~503_combout ;
wire \rfif.rdat1[6]~506_combout ;
wire \rfif.rdat1[6]~510_combout ;
wire \rfif.rdat1[6]~511_combout ;
wire \regs[2][6]~feeder_combout ;
wire \regs[2][6]~q ;
wire \rfif.rdat1[6]~515_combout ;
wire \regs[7][6]~feeder_combout ;
wire \regs[7][6]~q ;
wire \rfif.rdat1[6]~513_combout ;
wire \rfif.rdat1[6]~516_combout ;
wire \regs[13][6]~q ;
wire \regs[12][6]~q ;
wire \rfif.rdat1[6]~517_combout ;
wire \rfif.rdat1[6]~518_combout ;
wire \regs[28][5]~q ;
wire \regs[24][5]~q ;
wire \regs[16][5]~q ;
wire \rfif.rdat2[5]~550_combout ;
wire \rfif.rdat2[5]~551_combout ;
wire \rfif.rdat2[5]~552_combout ;
wire \regs[27][5]~q ;
wire \regs[31][5]~q ;
wire \rfif.rdat2[5]~554_combout ;
wire \regs[22][5]~q ;
wire \regs[30][5]~q ;
wire \rfif.rdat2[5]~547_combout ;
wire \rfif.rdat2[5]~555_combout ;
wire \regs[10][5]~q ;
wire \regs[11][5]~q ;
wire \regs[8][5]~q ;
wire \regs[9][5]~q ;
wire \rfif.rdat2[5]~556_combout ;
wire \rfif.rdat2[5]~557_combout ;
wire \regs[12][5]~feeder_combout ;
wire \regs[12][5]~q ;
wire \regs[14][5]~q ;
wire \rfif.rdat2[5]~563_combout ;
wire \regs[15][5]~q ;
wire \regs[13][5]~feeder_combout ;
wire \regs[13][5]~q ;
wire \rfif.rdat2[5]~564_combout ;
wire \regs[2][5]~q ;
wire \regs[3][5]~q ;
wire \regs[0][5]~q ;
wire \regs[1][5]~q ;
wire \rfif.rdat2[5]~560_combout ;
wire \rfif.rdat2[5]~561_combout ;
wire \regs[5][5]~q ;
wire \regs[7][5]~q ;
wire \regs[4][5]~q ;
wire \regs[6][5]~q ;
wire \rfif.rdat2[5]~558_combout ;
wire \rfif.rdat2[5]~559_combout ;
wire \rfif.rdat2[5]~562_combout ;
wire \rfif.rdat2[5]~565_combout ;
wire \regs[19][5]~q ;
wire \rfif.rdat1[5]~527_combout ;
wire \regs[23][5]~q ;
wire \rfif.rdat1[5]~528_combout ;
wire \regs[29][5]~q ;
wire \regs[21][5]~q ;
wire \regs[25][5]~q ;
wire \rfif.rdat1[5]~520_combout ;
wire \rfif.rdat1[5]~521_combout ;
wire \regs[26][5]~q ;
wire \rfif.rdat1[5]~523_combout ;
wire \rfif.rdat1[5]~525_combout ;
wire \rfif.rdat1[5]~526_combout ;
wire \rfif.rdat1[5]~530_combout ;
wire \rfif.rdat1[5]~531_combout ;
wire \rfif.rdat1[5]~537_combout ;
wire \rfif.rdat1[5]~538_combout ;
wire \rfif.rdat1[5]~534_combout ;
wire \rfif.rdat1[5]~535_combout ;
wire \rfif.rdat1[5]~532_combout ;
wire \rfif.rdat1[5]~533_combout ;
wire \rfif.rdat1[5]~536_combout ;
wire \regs[0][4]~q ;
wire \regs[2][4]~q ;
wire \rfif.rdat2[4]~581_combout ;
wire \regs[3][4]~q ;
wire \regs[1][4]~q ;
wire \rfif.rdat2[4]~582_combout ;
wire \rfif.rdat2[4]~583_combout ;
wire \regs[15][4]~q ;
wire \regs[14][4]~q ;
wire \regs[13][4]~q ;
wire \regs[12][4]~q ;
wire \rfif.rdat2[4]~584_combout ;
wire \rfif.rdat2[4]~585_combout ;
wire \regs[7][4]~feeder_combout ;
wire \regs[7][4]~q ;
wire \regs[6][4]~q ;
wire \regs[4][4]~q ;
wire \regs[5][4]~feeder_combout ;
wire \regs[5][4]~q ;
wire \rfif.rdat2[4]~577_combout ;
wire \rfif.rdat2[4]~578_combout ;
wire \rfif.rdat2[4]~586_combout ;
wire \regs[18][4]~q ;
wire \regs[22][4]~q ;
wire \rfif.rdat2[4]~569_combout ;
wire \regs[30][4]~q ;
wire \regs[26][4]~q ;
wire \rfif.rdat2[4]~570_combout ;
wire \regs[24][4]~q ;
wire \regs[28][4]~feeder_combout ;
wire \regs[28][4]~q ;
wire \regs[16][4]~q ;
wire \rfif.rdat2[4]~571_combout ;
wire \rfif.rdat2[4]~572_combout ;
wire \rfif.rdat2[4]~573_combout ;
wire \regs[21][4]~q ;
wire \regs[25][4]~q ;
wire \regs[17][4]~q ;
wire \rfif.rdat2[4]~567_combout ;
wire \rfif.rdat2[4]~568_combout ;
wire \regs[23][4]~q ;
wire \regs[31][4]~feeder_combout ;
wire \regs[31][4]~q ;
wire \rfif.rdat2[4]~575_combout ;
wire \rfif.rdat2[4]~576_combout ;
wire \regs[20][4]~feeder_combout ;
wire \regs[20][4]~q ;
wire \rfif.rdat1[4]~544_combout ;
wire \rfif.rdat1[4]~545_combout ;
wire \rfif.rdat1[4]~542_combout ;
wire \regs[29][4]~q ;
wire \rfif.rdat1[4]~543_combout ;
wire \rfif.rdat1[4]~546_combout ;
wire \regs[27][4]~q ;
wire \rfif.rdat1[4]~547_combout ;
wire \rfif.rdat1[4]~548_combout ;
wire \rfif.rdat1[4]~540_combout ;
wire \rfif.rdat1[4]~541_combout ;
wire \rfif.rdat1[4]~554_combout ;
wire \rfif.rdat1[4]~555_combout ;
wire \rfif.rdat1[4]~552_combout ;
wire \rfif.rdat1[4]~553_combout ;
wire \rfif.rdat1[4]~556_combout ;
wire \rfif.rdat1[4]~557_combout ;
wire \rfif.rdat1[4]~558_combout ;
wire \regs[11][4]~feeder_combout ;
wire \regs[11][4]~q ;
wire \regs[10][4]~feeder_combout ;
wire \regs[10][4]~q ;
wire \regs[9][4]~feeder_combout ;
wire \regs[9][4]~q ;
wire \regs[8][4]~feeder_combout ;
wire \regs[8][4]~q ;
wire \rfif.rdat1[4]~550_combout ;
wire \rfif.rdat1[4]~551_combout ;
wire \regs[22][3]~q ;
wire \regs[18][3]~q ;
wire \regs[26][3]~q ;
wire \rfif.rdat2[3]~588_combout ;
wire \rfif.rdat2[3]~589_combout ;
wire \regs[31][3]~q ;
wire \regs[27][3]~q ;
wire \rfif.rdat2[3]~596_combout ;
wire \regs[25][3]~q ;
wire \regs[29][3]~q ;
wire \regs[17][3]~q ;
wire \rfif.rdat2[3]~590_combout ;
wire \rfif.rdat2[3]~591_combout ;
wire \regs[28][3]~q ;
wire \regs[16][3]~q ;
wire \regs[24][3]~q ;
wire \rfif.rdat2[3]~592_combout ;
wire \rfif.rdat2[3]~593_combout ;
wire \rfif.rdat2[3]~594_combout ;
wire \rfif.rdat2[3]~597_combout ;
wire \regs[2][3]~q ;
wire \regs[3][3]~q ;
wire \rfif.rdat2[3]~603_combout ;
wire \rfif.rdat2[3]~604_combout ;
wire \regs[14][3]~q ;
wire \regs[12][3]~q ;
wire \rfif.rdat2[3]~605_combout ;
wire \regs[15][3]~q ;
wire \rfif.rdat2[3]~606_combout ;
wire \regs[10][3]~q ;
wire \regs[11][3]~q ;
wire \rfif.rdat2[3]~599_combout ;
wire \rfif.rdat2[3]~607_combout ;
wire \regs[23][3]~q ;
wire \regs[19][3]~q ;
wire \rfif.rdat1[3]~567_combout ;
wire \rfif.rdat1[3]~568_combout ;
wire \rfif.rdat1[3]~560_combout ;
wire \regs[21][3]~q ;
wire \rfif.rdat1[3]~561_combout ;
wire \regs[30][3]~q ;
wire \rfif.rdat1[3]~563_combout ;
wire \rfif.rdat1[3]~565_combout ;
wire \rfif.rdat1[3]~566_combout ;
wire \regs[5][3]~q ;
wire \rfif.rdat1[3]~570_combout ;
wire \regs[6][3]~q ;
wire \regs[7][3]~q ;
wire \rfif.rdat1[3]~571_combout ;
wire \rfif.rdat1[3]~574_combout ;
wire \regs[1][3]~q ;
wire \rfif.rdat1[3]~575_combout ;
wire \regs[9][3]~q ;
wire \regs[8][3]~q ;
wire \rfif.rdat1[3]~572_combout ;
wire \rfif.rdat1[3]~573_combout ;
wire \rfif.rdat1[3]~576_combout ;
wire \regs[13][3]~q ;
wire \rfif.rdat1[3]~577_combout ;
wire \rfif.rdat1[3]~578_combout ;
wire \regs[5][2]~q ;
wire \regs[4][2]~q ;
wire \rfif.rdat2[2]~619_combout ;
wire \regs[6][2]~q ;
wire \rfif.rdat2[2]~620_combout ;
wire \regs[8][2]~q ;
wire \regs[10][2]~q ;
wire \rfif.rdat2[2]~621_combout ;
wire \regs[11][2]~q ;
wire \regs[9][2]~q ;
wire \rfif.rdat2[2]~622_combout ;
wire \regs[2][2]~q ;
wire \regs[0][2]~q ;
wire \rfif.rdat2[2]~623_combout ;
wire \regs[3][2]~q ;
wire \regs[1][2]~feeder_combout ;
wire \regs[1][2]~q ;
wire \rfif.rdat2[2]~624_combout ;
wire \rfif.rdat2[2]~625_combout ;
wire \regs[12][2]~q ;
wire \regs[13][2]~q ;
wire \rfif.rdat2[2]~626_combout ;
wire \regs[15][2]~q ;
wire \regs[14][2]~q ;
wire \rfif.rdat2[2]~627_combout ;
wire \rfif.rdat2[2]~628_combout ;
wire \regs[23][2]~q ;
wire \regs[31][2]~q ;
wire \rfif.rdat2[2]~617_combout ;
wire \regs[29][2]~q ;
wire \regs[21][2]~q ;
wire \regs[17][2]~q ;
wire \regs[25][2]~q ;
wire \rfif.rdat2[2]~609_combout ;
wire \rfif.rdat2[2]~610_combout ;
wire \regs[16][2]~q ;
wire \regs[20][2]~q ;
wire \rfif.rdat2[2]~613_combout ;
wire \regs[28][2]~q ;
wire \regs[24][2]~q ;
wire \rfif.rdat2[2]~614_combout ;
wire \regs[26][2]~q ;
wire \regs[30][2]~q ;
wire \regs[18][2]~q ;
wire \regs[22][2]~q ;
wire \rfif.rdat2[2]~611_combout ;
wire \rfif.rdat2[2]~612_combout ;
wire \rfif.rdat2[2]~615_combout ;
wire \rfif.rdat2[2]~618_combout ;
wire \rfif.rdat1[2]~582_combout ;
wire \rfif.rdat1[2]~583_combout ;
wire \rfif.rdat1[2]~584_combout ;
wire \rfif.rdat1[2]~585_combout ;
wire \rfif.rdat1[2]~586_combout ;
wire \rfif.rdat1[2]~587_combout ;
wire \regs[27][2]~feeder_combout ;
wire \regs[27][2]~q ;
wire \rfif.rdat1[2]~588_combout ;
wire \rfif.rdat1[2]~580_combout ;
wire \rfif.rdat1[2]~581_combout ;
wire \rfif.rdat1[2]~597_combout ;
wire \rfif.rdat1[2]~598_combout ;
wire \rfif.rdat1[2]~590_combout ;
wire \rfif.rdat1[2]~591_combout ;
wire \rfif.rdat1[2]~594_combout ;
wire \rfif.rdat1[2]~595_combout ;
wire \rfif.rdat1[2]~592_combout ;
wire \regs[7][2]~q ;
wire \rfif.rdat1[2]~593_combout ;
wire \rfif.rdat1[2]~596_combout ;
wire \regs[27][1]~q ;
wire \regs[31][1]~q ;
wire \rfif.rdat2[1]~638_combout ;
wire \regs[22][1]~q ;
wire \regs[30][1]~q ;
wire \rfif.rdat2[1]~631_combout ;
wire \regs[28][1]~q ;
wire \regs[20][1]~q ;
wire \rfif.rdat2[1]~635_combout ;
wire \regs[17][1]~q ;
wire \regs[21][1]~q ;
wire \rfif.rdat2[1]~632_combout ;
wire \regs[29][1]~q ;
wire \regs[25][1]~q ;
wire \rfif.rdat2[1]~633_combout ;
wire \rfif.rdat2[1]~636_combout ;
wire \rfif.rdat2[1]~639_combout ;
wire \regs[13][1]~q ;
wire \regs[15][1]~q ;
wire \regs[14][1]~q ;
wire \regs[12][1]~q ;
wire \rfif.rdat2[1]~647_combout ;
wire \rfif.rdat2[1]~648_combout ;
wire \regs[5][1]~q ;
wire \regs[7][1]~q ;
wire \regs[6][1]~q ;
wire \regs[4][1]~q ;
wire \rfif.rdat2[1]~642_combout ;
wire \rfif.rdat2[1]~643_combout ;
wire \regs[2][1]~feeder_combout ;
wire \regs[2][1]~q ;
wire \regs[3][1]~q ;
wire \regs[0][1]~q ;
wire \regs[1][1]~q ;
wire \rfif.rdat2[1]~644_combout ;
wire \rfif.rdat2[1]~645_combout ;
wire \rfif.rdat2[1]~646_combout ;
wire \regs[10][1]~q ;
wire \regs[9][1]~q ;
wire \rfif.rdat2[1]~640_combout ;
wire \rfif.rdat2[1]~641_combout ;
wire \rfif.rdat2[1]~649_combout ;
wire \regs[26][1]~q ;
wire \regs[18][1]~q ;
wire \rfif.rdat1[1]~602_combout ;
wire \rfif.rdat1[1]~603_combout ;
wire \rfif.rdat1[1]~604_combout ;
wire \regs[24][1]~q ;
wire \rfif.rdat1[1]~605_combout ;
wire \rfif.rdat1[1]~606_combout ;
wire \regs[19][1]~q ;
wire \rfif.rdat1[1]~607_combout ;
wire \regs[23][1]~q ;
wire \rfif.rdat1[1]~608_combout ;
wire \rfif.rdat1[1]~600_combout ;
wire \rfif.rdat1[1]~601_combout ;
wire \rfif.rdat1[1]~614_combout ;
wire \rfif.rdat1[1]~615_combout ;
wire \regs[11][1]~q ;
wire \regs[8][1]~q ;
wire \rfif.rdat1[1]~612_combout ;
wire \rfif.rdat1[1]~613_combout ;
wire \rfif.rdat1[1]~616_combout ;
wire \rfif.rdat1[1]~617_combout ;
wire \rfif.rdat1[1]~618_combout ;
wire \rfif.rdat1[1]~610_combout ;
wire \rfif.rdat1[1]~611_combout ;
wire \regs[0][0]~q ;
wire \regs[2][0]~q ;
wire \rfif.rdat2[0]~665_combout ;
wire \regs[3][0]~q ;
wire \regs[1][0]~q ;
wire \rfif.rdat2[0]~666_combout ;
wire \rfif.rdat2[0]~667_combout ;
wire \regs[12][0]~q ;
wire \regs[13][0]~q ;
wire \rfif.rdat2[0]~668_combout ;
wire \regs[15][0]~feeder_combout ;
wire \regs[15][0]~q ;
wire \rfif.rdat2[0]~669_combout ;
wire \regs[6][0]~q ;
wire \regs[7][0]~q ;
wire \rfif.rdat2[0]~662_combout ;
wire \rfif.rdat2[0]~670_combout ;
wire \regs[28][0]~q ;
wire \regs[24][0]~q ;
wire \rfif.rdat2[0]~656_combout ;
wire \regs[30][0]~q ;
wire \regs[26][0]~q ;
wire \rfif.rdat2[0]~654_combout ;
wire \rfif.rdat2[0]~657_combout ;
wire \regs[17][0]~q ;
wire \regs[25][0]~q ;
wire \rfif.rdat2[0]~651_combout ;
wire \regs[21][0]~q ;
wire \regs[29][0]~q ;
wire \rfif.rdat2[0]~652_combout ;
wire \regs[23][0]~q ;
wire \regs[31][0]~q ;
wire \rfif.rdat2[0]~659_combout ;
wire \rfif.rdat2[0]~660_combout ;
wire \regs[22][0]~q ;
wire \regs[18][0]~q ;
wire \rfif.rdat1[0]~620_combout ;
wire \rfif.rdat1[0]~621_combout ;
wire \rfif.rdat1[0]~627_combout ;
wire \regs[27][0]~q ;
wire \rfif.rdat1[0]~628_combout ;
wire \rfif.rdat1[0]~622_combout ;
wire \rfif.rdat1[0]~623_combout ;
wire \rfif.rdat1[0]~624_combout ;
wire \regs[20][0]~q ;
wire \rfif.rdat1[0]~625_combout ;
wire \rfif.rdat1[0]~626_combout ;
wire \regs[8][0]~q ;
wire \regs[9][0]~q ;
wire \rfif.rdat1[0]~630_combout ;
wire \regs[10][0]~q ;
wire \regs[11][0]~q ;
wire \rfif.rdat1[0]~631_combout ;
wire \regs[14][0]~q ;
wire \rfif.rdat1[0]~637_combout ;
wire \rfif.rdat1[0]~638_combout ;
wire \rfif.rdat1[0]~634_combout ;
wire \rfif.rdat1[0]~635_combout ;
wire \regs[5][0]~q ;
wire \regs[4][0]~q ;
wire \rfif.rdat1[0]~632_combout ;
wire \rfif.rdat1[0]~633_combout ;
wire \rfif.rdat1[0]~636_combout ;


// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[31]~2 (
// Equation(s):
// \rfif.rdat2[31]~2_combout  = (Instr_IF_18 & ((\regs[21][31]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[17][31]~q  & !Instr_IF_19))))

	.dataa(Instr_IF_18),
	.datab(\regs[21][31]~q ),
	.datac(\regs[17][31]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~2_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~2 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[31]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \regs[29][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][31] .is_wysiwyg = "true";
defparam \regs[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[31]~3 (
// Equation(s):
// \rfif.rdat2[31]~3_combout  = (Instr_IF_19 & ((\rfif.rdat2[31]~2_combout  & (\regs[29][31]~q )) # (!\rfif.rdat2[31]~2_combout  & ((\regs[25][31]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[31]~2_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[31]~2_combout ),
	.datac(\regs[29][31]~q ),
	.datad(\regs[25][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~3 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N13
dffeas \regs[20][31] (
	.clk(!CLK),
	.d(\regs[20][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][31] .is_wysiwyg = "true";
defparam \regs[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[31]~7 (
// Equation(s):
// \rfif.rdat2[31]~7_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[23][31]~q )) # (!Instr_IF_18 & ((\regs[19][31]~q )))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[23][31]~q ),
	.datad(\regs[19][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~7_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~7 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[31]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N12
cycloneive_lcell_comb \rfif.rdat2[31]~10 (
// Equation(s):
// \rfif.rdat2[31]~10_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[9][31]~q ))) # (!Instr_IF_16 & (\regs[8][31]~q ))))

	.dataa(Instr_IF_17),
	.datab(\regs[8][31]~q ),
	.datac(\regs[9][31]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~10_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~10 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[31]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N13
dffeas \regs[1][31] (
	.clk(!CLK),
	.d(\regs[1][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][31] .is_wysiwyg = "true";
defparam \regs[1][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N15
dffeas \regs[0][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][31] .is_wysiwyg = "true";
defparam \regs[0][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[31]~14 (
// Equation(s):
// \rfif.rdat2[31]~14_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[1][31]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[0][31]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][31]~q ),
	.datad(\regs[1][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~14_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~14 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[31]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \rfif.rdat2[31]~15 (
// Equation(s):
// \rfif.rdat2[31]~15_combout  = (Instr_IF_17 & ((\rfif.rdat2[31]~14_combout  & ((\regs[3][31]~q ))) # (!\rfif.rdat2[31]~14_combout  & (\regs[2][31]~q )))) # (!Instr_IF_17 & (\rfif.rdat2[31]~14_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[31]~14_combout ),
	.datac(\regs[2][31]~q ),
	.datad(\regs[3][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~15_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~15 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[31]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[31]~17 (
// Equation(s):
// \rfif.rdat2[31]~17_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][31]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][31]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][31]~q ),
	.datad(\regs[14][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~17_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~17 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[31]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[31]~14 (
// Equation(s):
// \rfif.rdat1[31]~14_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][31]~q )) # (!Instr_IF_21 & ((\regs[0][31]~q )))))

	.dataa(Instr_IF_22),
	.datab(\regs[1][31]~q ),
	.datac(Instr_IF_21),
	.datad(\regs[0][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~14_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~14 .lut_mask = 16'hE5E0;
defparam \rfif.rdat1[31]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N15
dffeas \regs[19][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][30] .is_wysiwyg = "true";
defparam \regs[19][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \regs[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][30] .is_wysiwyg = "true";
defparam \regs[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \rfif.rdat2[30]~28 (
// Equation(s):
// \rfif.rdat2[30]~28_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\regs[27][30]~q )) # (!Instr_IF_19 & ((\regs[19][30]~q )))))

	.dataa(Instr_IF_18),
	.datab(\regs[27][30]~q ),
	.datac(\regs[19][30]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~28_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~28 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[30]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \rfif.rdat2[30]~38 (
// Equation(s):
// \rfif.rdat2[30]~38_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][30]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][30]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][30]~q ),
	.datad(\regs[13][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~38_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~38 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[30]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N21
dffeas \regs[21][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][29] .is_wysiwyg = "true";
defparam \regs[21][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N7
dffeas \regs[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][29] .is_wysiwyg = "true";
defparam \regs[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[29]~42 (
// Equation(s):
// \rfif.rdat1[29]~42_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[21][29]~q )) # (!Instr_IF_23 & ((\regs[17][29]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[21][29]~q ),
	.datad(\regs[17][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~42_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~42 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[29]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N23
dffeas \regs[28][29] (
	.clk(!CLK),
	.d(\regs[28][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][29] .is_wysiwyg = "true";
defparam \regs[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N27
dffeas \regs[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][29] .is_wysiwyg = "true";
defparam \regs[3][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N31
dffeas \regs[12][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][29] .is_wysiwyg = "true";
defparam \regs[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[29]~44 (
// Equation(s):
// \rfif.rdat2[29]~44_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[21][29]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[17][29]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][29]~q ),
	.datad(\regs[21][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~44_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~44 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[29]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N24
cycloneive_lcell_comb \rfif.rdat2[29]~46 (
// Equation(s):
// \rfif.rdat2[29]~46_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[24][29]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[16][29]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][29]~q ),
	.datad(\regs[24][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~46_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~46 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[29]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[29]~47 (
// Equation(s):
// \rfif.rdat2[29]~47_combout  = (Instr_IF_18 & ((\rfif.rdat2[29]~46_combout  & (\regs[28][29]~q )) # (!\rfif.rdat2[29]~46_combout  & ((\regs[20][29]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[29]~46_combout ))))

	.dataa(\regs[28][29]~q ),
	.datab(\regs[20][29]~q ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[29]~46_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~47_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~47 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[29]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \rfif.rdat2[29]~56 (
// Equation(s):
// \rfif.rdat2[29]~56_combout  = (Instr_IF_16 & ((\regs[1][29]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((!Instr_IF_17 & \regs[0][29]~q ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][29]~q ),
	.datac(Instr_IF_17),
	.datad(\regs[0][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~56_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~56 .lut_mask = 16'hADA8;
defparam \rfif.rdat2[29]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[29]~57 (
// Equation(s):
// \rfif.rdat2[29]~57_combout  = (Instr_IF_17 & ((\rfif.rdat2[29]~56_combout  & (\regs[3][29]~q )) # (!\rfif.rdat2[29]~56_combout  & ((\regs[2][29]~q ))))) # (!Instr_IF_17 & (\rfif.rdat2[29]~56_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[29]~56_combout ),
	.datac(\regs[3][29]~q ),
	.datad(\regs[2][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~57_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~57 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[29]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \rfif.rdat2[29]~59 (
// Equation(s):
// \rfif.rdat2[29]~59_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[14][29]~q ))) # (!Instr_IF_17 & (\regs[12][29]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][29]~q ),
	.datad(\regs[14][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~59_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~59 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[29]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N28
cycloneive_lcell_comb \rfif.rdat1[28]~72 (
// Equation(s):
// \rfif.rdat1[28]~72_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[10][28]~q ))) # (!Instr_IF_22 & (\regs[8][28]~q ))))

	.dataa(\regs[8][28]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[10][28]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~72_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~72 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[28]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N23
dffeas \regs[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][27] .is_wysiwyg = "true";
defparam \regs[6][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \rfif.rdat1[27]~92 (
// Equation(s):
// \rfif.rdat1[27]~92_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][27]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][27]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][27]~q ),
	.datad(\regs[4][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~92_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~92 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[27]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N27
dffeas \regs[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][26] .is_wysiwyg = "true";
defparam \regs[18][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N7
dffeas \regs[3][26] (
	.clk(!CLK),
	.d(\regs[3][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][26] .is_wysiwyg = "true";
defparam \regs[3][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[26]~105 (
// Equation(s):
// \rfif.rdat2[26]~105_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\regs[25][26]~q )) # (!Instr_IF_19 & ((\regs[17][26]~q )))))

	.dataa(Instr_IF_18),
	.datab(\regs[25][26]~q ),
	.datac(\regs[17][26]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~105_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~105 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[26]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \rfif.rdat2[26]~107 (
// Equation(s):
// \rfif.rdat2[26]~107_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[22][26]~q )) # (!Instr_IF_18 & ((\regs[18][26]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[22][26]~q ),
	.datac(\regs[18][26]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~107_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~107 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[26]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[26]~108 (
// Equation(s):
// \rfif.rdat2[26]~108_combout  = (Instr_IF_19 & ((\rfif.rdat2[26]~107_combout  & ((\regs[30][26]~q ))) # (!\rfif.rdat2[26]~107_combout  & (\regs[26][26]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[26]~107_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][26]~q ),
	.datac(\regs[30][26]~q ),
	.datad(\rfif.rdat2[26]~107_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~108_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~108 .lut_mask = 16'hF588;
defparam \rfif.rdat2[26]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \rfif.rdat2[26]~122 (
// Equation(s):
// \rfif.rdat2[26]~122_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][26]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][26]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][26]~q ),
	.datad(\regs[13][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~122_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~122 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[26]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[25]~122 (
// Equation(s):
// \rfif.rdat1[25]~122_combout  = (Instr_IF_23 & (((\regs[21][25]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[17][25]~q  & ((!Instr_IF_24))))

	.dataa(\regs[17][25]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[21][25]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~122_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~122 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[25]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N7
dffeas \regs[28][25] (
	.clk(!CLK),
	.d(\regs[28][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][25] .is_wysiwyg = "true";
defparam \regs[28][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[25]~132 (
// Equation(s):
// \rfif.rdat1[25]~132_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][25]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][25]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][25]~q ),
	.datad(\regs[4][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~132_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~132 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[25]~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \rfif.rdat2[25]~140 (
// Equation(s):
// \rfif.rdat2[25]~140_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[1][25]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[0][25]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][25]~q ),
	.datad(\regs[1][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~140_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~140 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[25]~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[25]~141 (
// Equation(s):
// \rfif.rdat2[25]~141_combout  = (Instr_IF_17 & ((\rfif.rdat2[25]~140_combout  & (\regs[3][25]~q )) # (!\rfif.rdat2[25]~140_combout  & ((\regs[2][25]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[25]~140_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[3][25]~q ),
	.datac(\regs[2][25]~q ),
	.datad(\rfif.rdat2[25]~140_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~141_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~141 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[25]~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N11
dffeas \regs[28][24] (
	.clk(!CLK),
	.d(\regs[28][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][24] .is_wysiwyg = "true";
defparam \regs[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N31
dffeas \regs[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][24] .is_wysiwyg = "true";
defparam \regs[8][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N11
dffeas \regs[3][24] (
	.clk(!CLK),
	.d(\regs[3][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][24] .is_wysiwyg = "true";
defparam \regs[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[24]~151 (
// Equation(s):
// \rfif.rdat2[24]~151_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][24]~q ))) # (!Instr_IF_18 & (\regs[16][24]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][24]~q ),
	.datad(\regs[20][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~151_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~151 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[24]~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[24]~152 (
// Equation(s):
// \rfif.rdat2[24]~152_combout  = (\rfif.rdat2[24]~151_combout  & ((\regs[28][24]~q ) # ((!Instr_IF_19)))) # (!\rfif.rdat2[24]~151_combout  & (((\regs[24][24]~q  & Instr_IF_19))))

	.dataa(\regs[28][24]~q ),
	.datab(\regs[24][24]~q ),
	.datac(\rfif.rdat2[24]~151_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~152_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~152 .lut_mask = 16'hACF0;
defparam \rfif.rdat2[24]~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[24]~154 (
// Equation(s):
// \rfif.rdat2[24]~154_combout  = (Instr_IF_19 & ((\regs[27][24]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[19][24]~q  & !Instr_IF_18))))

	.dataa(\regs[27][24]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[19][24]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~154_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~154 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[24]~154 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[24]~159 (
// Equation(s):
// \rfif.rdat2[24]~159_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][24]~q ))) # (!Instr_IF_17 & (\regs[8][24]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][24]~q ),
	.datad(\regs[10][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~159_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~159 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[24]~159 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[24]~160 (
// Equation(s):
// \rfif.rdat2[24]~160_combout  = (Instr_IF_16 & ((\rfif.rdat2[24]~159_combout  & (\regs[11][24]~q )) # (!\rfif.rdat2[24]~159_combout  & ((\regs[9][24]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[24]~159_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[24]~159_combout ),
	.datac(\regs[11][24]~q ),
	.datad(\regs[9][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~160_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~160 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[24]~160 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N31
dffeas \regs[28][23] (
	.clk(!CLK),
	.d(\regs[28][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][23] .is_wysiwyg = "true";
defparam \regs[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N31
dffeas \regs[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][23] .is_wysiwyg = "true";
defparam \regs[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \rfif.rdat2[23]~168 (
// Equation(s):
// \rfif.rdat2[23]~168_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][23]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][23]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][23]~q ),
	.datad(\regs[26][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~168_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~168 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[23]~168 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \rfif.rdat2[23]~178 (
// Equation(s):
// \rfif.rdat2[23]~178_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][23]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][23]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][23]~q ),
	.datad(\regs[9][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~178_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~178 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[23]~178 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[23]~180 (
// Equation(s):
// \rfif.rdat2[23]~180_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][23]~q ))) # (!Instr_IF_17 & (\regs[4][23]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][23]~q ),
	.datad(\regs[6][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~180_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~180 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[23]~180 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[22]~184 (
// Equation(s):
// \rfif.rdat1[22]~184_combout  = (Instr_IF_23 & (((\regs[20][22]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][22]~q  & ((!Instr_IF_24))))

	.dataa(\regs[16][22]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][22]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~184_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~184 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[22]~184 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N13
dffeas \regs[1][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][22] .is_wysiwyg = "true";
defparam \regs[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[22]~199 (
// Equation(s):
// \rfif.rdat2[22]~199_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][22]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][22]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][22]~q ),
	.datad(\regs[5][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~199_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~199 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[22]~199 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \rfif.rdat2[22]~201 (
// Equation(s):
// \rfif.rdat2[22]~201_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][22]~q ))) # (!Instr_IF_17 & (\regs[8][22]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][22]~q ),
	.datad(\regs[10][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~201_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~201 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[22]~201 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \rfif.rdat2[22]~206 (
// Equation(s):
// \rfif.rdat2[22]~206_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[13][22]~q ))) # (!Instr_IF_16 & (\regs[12][22]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][22]~q ),
	.datad(\regs[13][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~206_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~206 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[22]~206 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N29
dffeas \regs[24][21] (
	.clk(!CLK),
	.d(\regs[24][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][21] .is_wysiwyg = "true";
defparam \regs[24][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \regs[16][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][21] .is_wysiwyg = "true";
defparam \regs[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[21]~204 (
// Equation(s):
// \rfif.rdat1[21]~204_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][21]~q ))) # (!Instr_IF_24 & (\regs[16][21]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[16][21]~q ),
	.datad(\regs[24][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~204_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~204 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[21]~204 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \rfif.rdat1[21]~214 (
// Equation(s):
// \rfif.rdat1[21]~214_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[1][21]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & (\regs[0][21]~q )))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[0][21]~q ),
	.datad(\regs[1][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~214_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~214 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[21]~214 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \rfif.rdat2[21]~214 (
// Equation(s):
// \rfif.rdat2[21]~214_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][21]~q ))) # (!Instr_IF_19 & (\regs[16][21]~q ))))

	.dataa(\regs[16][21]~q ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\regs[24][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~214_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~214 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[21]~214 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[21]~215 (
// Equation(s):
// \rfif.rdat2[21]~215_combout  = (Instr_IF_18 & ((\rfif.rdat2[21]~214_combout  & (\regs[28][21]~q )) # (!\rfif.rdat2[21]~214_combout  & ((\regs[20][21]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[21]~214_combout ))))

	.dataa(\regs[28][21]~q ),
	.datab(\regs[20][21]~q ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[21]~214_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~215_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~215 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[21]~215 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \rfif.rdat2[21]~220 (
// Equation(s):
// \rfif.rdat2[21]~220_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[9][21]~q ))) # (!Instr_IF_16 & (\regs[8][21]~q ))))

	.dataa(\regs[8][21]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[9][21]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~220_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~220 .lut_mask = 16'hFC22;
defparam \rfif.rdat2[21]~220 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \rfif.rdat2[21]~222 (
// Equation(s):
// \rfif.rdat2[21]~222_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][21]~q ))) # (!Instr_IF_17 & (\regs[4][21]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][21]~q ),
	.datad(\regs[6][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~222_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~222 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[21]~222 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \rfif.rdat2[21]~223 (
// Equation(s):
// \rfif.rdat2[21]~223_combout  = (Instr_IF_16 & ((\rfif.rdat2[21]~222_combout  & (\regs[7][21]~q )) # (!\rfif.rdat2[21]~222_combout  & ((\regs[5][21]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[21]~222_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[7][21]~q ),
	.datac(\rfif.rdat2[21]~222_combout ),
	.datad(\regs[5][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~223_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~223 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[21]~223 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N7
dffeas \regs[16][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][20] .is_wysiwyg = "true";
defparam \regs[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[20]~235 (
// Equation(s):
// \rfif.rdat2[20]~235_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[20][20]~q )) # (!Instr_IF_18 & ((\regs[16][20]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[20][20]~q ),
	.datac(\regs[16][20]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~235_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~235 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[20]~235 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[19]~242 (
// Equation(s):
// \rfif.rdat1[19]~242_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][19]~q ))) # (!Instr_IF_23 & (\regs[17][19]~q ))))

	.dataa(\regs[17][19]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[21][19]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~242_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~242 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[19]~242 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \rfif.rdat1[19]~244 (
// Equation(s):
// \rfif.rdat1[19]~244_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[24][19]~q )) # (!Instr_IF_24 & ((\regs[16][19]~q )))))

	.dataa(\regs[24][19]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[16][19]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~244_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~244 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[19]~244 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \rfif.rdat1[19]~252 (
// Equation(s):
// \rfif.rdat1[19]~252_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[6][19]~q ))) # (!Instr_IF_22 & (\regs[4][19]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[4][19]~q ),
	.datac(\regs[6][19]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~252_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~252 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[19]~252 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N5
dffeas \regs[2][19] (
	.clk(!CLK),
	.d(\regs[2][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][19] .is_wysiwyg = "true";
defparam \regs[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N13
dffeas \regs[1][19] (
	.clk(!CLK),
	.d(\regs[1][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][19] .is_wysiwyg = "true";
defparam \regs[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \rfif.rdat2[19]~269 (
// Equation(s):
// \rfif.rdat2[19]~269_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][19]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][19]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][19]~q ),
	.datad(\regs[14][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~269_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~269 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[19]~269 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[18]~273 (
// Equation(s):
// \rfif.rdat2[18]~273_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[25][18]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[17][18]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][18]~q ),
	.datad(\regs[25][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~273_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~273 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[18]~273 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N27
dffeas \regs[16][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][17] .is_wysiwyg = "true";
defparam \regs[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[17]~284 (
// Equation(s):
// \rfif.rdat1[17]~284_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[24][17]~q )) # (!Instr_IF_24 & ((\regs[16][17]~q )))))

	.dataa(\regs[24][17]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[16][17]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~284_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~284 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[17]~284 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[17]~292 (
// Equation(s):
// \rfif.rdat1[17]~292_combout  = (Instr_IF_22 & (((Instr_IF_21) # (\regs[6][17]~q )))) # (!Instr_IF_22 & (\regs[4][17]~q  & (!Instr_IF_21)))

	.dataa(Instr_IF_22),
	.datab(\regs[4][17]~q ),
	.datac(Instr_IF_21),
	.datad(\regs[6][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~292_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~292 .lut_mask = 16'hAEA4;
defparam \rfif.rdat1[17]~292 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N15
dffeas \regs[2][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][17] .is_wysiwyg = "true";
defparam \regs[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \rfif.rdat2[17]~308 (
// Equation(s):
// \rfif.rdat2[17]~308_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][17]~q ))) # (!Instr_IF_16 & (\regs[0][17]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][17]~q ),
	.datad(\regs[1][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~308_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~308 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[17]~308 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[17]~309 (
// Equation(s):
// \rfif.rdat2[17]~309_combout  = (Instr_IF_17 & ((\rfif.rdat2[17]~308_combout  & ((\regs[3][17]~q ))) # (!\rfif.rdat2[17]~308_combout  & (\regs[2][17]~q )))) # (!Instr_IF_17 & (\rfif.rdat2[17]~308_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[17]~308_combout ),
	.datac(\regs[2][17]~q ),
	.datad(\regs[3][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~309_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~309 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[17]~309 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N21
dffeas \regs[22][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][16] .is_wysiwyg = "true";
defparam \regs[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N7
dffeas \regs[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][16] .is_wysiwyg = "true";
defparam \regs[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \rfif.rdat1[16]~302 (
// Equation(s):
// \rfif.rdat1[16]~302_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[22][16]~q )) # (!Instr_IF_23 & ((\regs[18][16]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[22][16]~q ),
	.datad(\regs[18][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~302_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~302 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[16]~302 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N25
dffeas \regs[20][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][16] .is_wysiwyg = "true";
defparam \regs[20][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N15
dffeas \regs[16][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][16] .is_wysiwyg = "true";
defparam \regs[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[16]~304 (
// Equation(s):
// \rfif.rdat1[16]~304_combout  = (Instr_IF_23 & (((\regs[20][16]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][16]~q  & ((!Instr_IF_24))))

	.dataa(\regs[16][16]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][16]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~304_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~304 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[16]~304 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N27
dffeas \regs[3][16] (
	.clk(!CLK),
	.d(\regs[3][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][16] .is_wysiwyg = "true";
defparam \regs[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \rfif.rdat2[16]~317 (
// Equation(s):
// \rfif.rdat2[16]~317_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][16]~q ))) # (!Instr_IF_18 & (\regs[18][16]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][16]~q ),
	.datad(\regs[22][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~317_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~317 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[16]~317 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \rfif.rdat2[16]~318 (
// Equation(s):
// \rfif.rdat2[16]~318_combout  = (\rfif.rdat2[16]~317_combout  & (((\regs[30][16]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[16]~317_combout  & (\regs[26][16]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[16]~317_combout ),
	.datab(\regs[26][16]~q ),
	.datac(\regs[30][16]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~318_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~318 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[16]~318 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[16]~319 (
// Equation(s):
// \rfif.rdat2[16]~319_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][16]~q ))) # (!Instr_IF_18 & (\regs[16][16]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][16]~q ),
	.datad(\regs[20][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~319_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~319 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[16]~319 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \rfif.rdat2[16]~327 (
// Equation(s):
// \rfif.rdat2[16]~327_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][16]~q ))) # (!Instr_IF_17 & (\regs[8][16]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][16]~q ),
	.datad(\regs[10][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~327_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~327 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[16]~327 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[15]~332 (
// Equation(s):
// \rfif.rdat1[15]~332_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][15]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][15]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][15]~q ),
	.datad(\regs[4][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~332_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~332 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[15]~332 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \rfif.rdat2[15]~343 (
// Equation(s):
// \rfif.rdat2[15]~343_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[23][15]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[19][15]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][15]~q ),
	.datad(\regs[23][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~343_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~343 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[15]~343 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N11
dffeas \regs[16][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][14] .is_wysiwyg = "true";
defparam \regs[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N10
cycloneive_lcell_comb \rfif.rdat1[14]~344 (
// Equation(s):
// \rfif.rdat1[14]~344_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[20][14]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[16][14]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[16][14]~q ),
	.datad(\regs[20][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~344_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~344 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[14]~344 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[14]~357 (
// Equation(s):
// \rfif.rdat2[14]~357_combout  = (Instr_IF_19 & ((\regs[25][14]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[17][14]~q  & !Instr_IF_18))))

	.dataa(\regs[25][14]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[17][14]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~357_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~357 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[14]~357 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N1
dffeas \regs[20][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][13] .is_wysiwyg = "true";
defparam \regs[20][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N27
dffeas \regs[16][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][13] .is_wysiwyg = "true";
defparam \regs[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[13]~382 (
// Equation(s):
// \rfif.rdat2[13]~382_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][13]~q ))) # (!Instr_IF_19 & (\regs[16][13]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][13]~q ),
	.datad(\regs[24][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~382_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~382 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[13]~382 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N30
cycloneive_lcell_comb \rfif.rdat2[13]~383 (
// Equation(s):
// \rfif.rdat2[13]~383_combout  = (Instr_IF_18 & ((\rfif.rdat2[13]~382_combout  & ((\regs[28][13]~q ))) # (!\rfif.rdat2[13]~382_combout  & (\regs[20][13]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[13]~382_combout ))))

	.dataa(\regs[20][13]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][13]~q ),
	.datad(\rfif.rdat2[13]~382_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~383_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~383 .lut_mask = 16'hF388;
defparam \rfif.rdat2[13]~383 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N13
dffeas \regs[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][13] .is_wysiwyg = "true";
defparam \regs[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[13]~390 (
// Equation(s):
// \rfif.rdat2[13]~390_combout  = (Instr_IF_17 & ((\regs[6][13]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\regs[4][13]~q  & !Instr_IF_16))))

	.dataa(\regs[6][13]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[4][13]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~390_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~390 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[13]~390 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[13]~391 (
// Equation(s):
// \rfif.rdat2[13]~391_combout  = (\rfif.rdat2[13]~390_combout  & ((\regs[7][13]~q ) # ((!Instr_IF_16)))) # (!\rfif.rdat2[13]~390_combout  & (((Instr_IF_16 & \regs[5][13]~q ))))

	.dataa(\rfif.rdat2[13]~390_combout ),
	.datab(\regs[7][13]~q ),
	.datac(Instr_IF_16),
	.datad(\regs[5][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~391_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~391 .lut_mask = 16'hDA8A;
defparam \rfif.rdat2[13]~391 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[13]~364 (
// Equation(s):
// \rfif.rdat1[13]~364_combout  = (Instr_IF_23 & (((\regs[20][13]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][13]~q  & ((!Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][13]~q ),
	.datac(\regs[20][13]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~364_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~364 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[13]~364 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N9
dffeas \regs[19][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][12] .is_wysiwyg = "true";
defparam \regs[19][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[12]~406 (
// Equation(s):
// \rfif.rdat2[12]~406_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[27][12]~q ))) # (!Instr_IF_19 & (\regs[19][12]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][12]~q ),
	.datad(\regs[27][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~406_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~406 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[12]~406 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N11
dffeas \regs[7][12] (
	.clk(!CLK),
	.d(\regs[7][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][12] .is_wysiwyg = "true";
defparam \regs[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \rfif.rdat2[12]~416 (
// Equation(s):
// \rfif.rdat2[12]~416_combout  = (Instr_IF_16 & ((\regs[13][12]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[12][12]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[13][12]~q ),
	.datac(\regs[12][12]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~416_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~416 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[12]~416 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[12]~394 (
// Equation(s):
// \rfif.rdat1[12]~394_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[1][12]~q ))) # (!Instr_IF_21 & (\regs[0][12]~q ))))

	.dataa(\regs[0][12]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[1][12]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~394_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~394 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[12]~394 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N7
dffeas \regs[16][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][11] .is_wysiwyg = "true";
defparam \regs[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[11]~424 (
// Equation(s):
// \rfif.rdat2[11]~424_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][11]~q ))) # (!Instr_IF_19 & (\regs[16][11]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][11]~q ),
	.datad(\regs[24][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~424_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~424 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[11]~424 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[11]~434 (
// Equation(s):
// \rfif.rdat2[11]~434_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][11]~q ))) # (!Instr_IF_16 & (\regs[0][11]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][11]~q ),
	.datad(\regs[1][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~434_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~434 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[11]~434 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[11]~435 (
// Equation(s):
// \rfif.rdat2[11]~435_combout  = (Instr_IF_17 & ((\rfif.rdat2[11]~434_combout  & ((\regs[3][11]~q ))) # (!\rfif.rdat2[11]~434_combout  & (\regs[2][11]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[11]~434_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[2][11]~q ),
	.datac(\regs[3][11]~q ),
	.datad(\rfif.rdat2[11]~434_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~435_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~435 .lut_mask = 16'hF588;
defparam \rfif.rdat2[11]~435 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N11
dffeas \regs[1][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][10] .is_wysiwyg = "true";
defparam \regs[1][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N7
dffeas \regs[0][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][10] .is_wysiwyg = "true";
defparam \regs[0][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[10]~455 (
// Equation(s):
// \rfif.rdat2[10]~455_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][10]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][10]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][10]~q ),
	.datad(\regs[2][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~455_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~455 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[10]~455 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[10]~456 (
// Equation(s):
// \rfif.rdat2[10]~456_combout  = (Instr_IF_16 & ((\rfif.rdat2[10]~455_combout  & ((\regs[3][10]~q ))) # (!\rfif.rdat2[10]~455_combout  & (\regs[1][10]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[10]~455_combout ))))

	.dataa(\regs[1][10]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[3][10]~q ),
	.datad(\rfif.rdat2[10]~455_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~456_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~456 .lut_mask = 16'hF388;
defparam \rfif.rdat2[10]~456 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \rfif.rdat1[10]~432 (
// Equation(s):
// \rfif.rdat1[10]~432_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][10]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][10]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][10]~q ),
	.datad(\regs[4][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~432_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~432 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[10]~432 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[10]~434 (
// Equation(s):
// \rfif.rdat1[10]~434_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][10]~q )) # (!Instr_IF_21 & ((\regs[0][10]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][10]~q ),
	.datad(\regs[0][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~434_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~434 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[10]~434 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \rfif.rdat2[9]~462 (
// Equation(s):
// \rfif.rdat2[9]~462_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[26][9]~q ))) # (!Instr_IF_19 & (\regs[18][9]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[18][9]~q ),
	.datac(\regs[26][9]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~462_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~462 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[9]~462 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[9]~464 (
// Equation(s):
// \rfif.rdat2[9]~464_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][9]~q ))) # (!Instr_IF_18 & (\regs[17][9]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][9]~q ),
	.datad(\regs[21][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~464_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~464 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[9]~464 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N17
dffeas \regs[20][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][9] .is_wysiwyg = "true";
defparam \regs[20][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N7
dffeas \regs[9][9] (
	.clk(!CLK),
	.d(\regs[9][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][9] .is_wysiwyg = "true";
defparam \regs[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N27
dffeas \regs[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][9] .is_wysiwyg = "true";
defparam \regs[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[9]~472 (
// Equation(s):
// \rfif.rdat2[9]~472_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][9]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][9]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][9]~q ),
	.datad(\regs[9][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~472_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~472 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[9]~472 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[9]~444 (
// Equation(s):
// \rfif.rdat1[9]~444_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[20][9]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & ((\regs[16][9]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[20][9]~q ),
	.datad(\regs[16][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~444_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~444 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[9]~444 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[9]~454 (
// Equation(s):
// \rfif.rdat1[9]~454_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][9]~q )) # (!Instr_IF_22 & ((\regs[0][9]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[2][9]~q ),
	.datad(\regs[0][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~454_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~454 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[9]~454 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \rfif.rdat2[8]~485 (
// Equation(s):
// \rfif.rdat2[8]~485_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][8]~q ))) # (!Instr_IF_18 & (\regs[18][8]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][8]~q ),
	.datad(\regs[22][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~485_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~485 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[8]~485 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N5
dffeas \regs[24][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][8] .is_wysiwyg = "true";
defparam \regs[24][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N3
dffeas \regs[16][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][8] .is_wysiwyg = "true";
defparam \regs[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N2
cycloneive_lcell_comb \rfif.rdat2[8]~487 (
// Equation(s):
// \rfif.rdat2[8]~487_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[20][8]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[16][8]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][8]~q ),
	.datad(\regs[20][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~487_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~487 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[8]~487 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \rfif.rdat2[8]~488 (
// Equation(s):
// \rfif.rdat2[8]~488_combout  = (Instr_IF_19 & ((\rfif.rdat2[8]~487_combout  & ((\regs[28][8]~q ))) # (!\rfif.rdat2[8]~487_combout  & (\regs[24][8]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[8]~487_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[24][8]~q ),
	.datac(\regs[28][8]~q ),
	.datad(\rfif.rdat2[8]~487_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~488_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~488 .lut_mask = 16'hF588;
defparam \rfif.rdat2[8]~488 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[8]~464 (
// Equation(s):
// \rfif.rdat1[8]~464_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][8]~q ))) # (!Instr_IF_24 & (\regs[16][8]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][8]~q ),
	.datac(\regs[24][8]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~464_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~464 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[8]~464 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N19
dffeas \regs[16][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][7] .is_wysiwyg = "true";
defparam \regs[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[7]~508 (
// Equation(s):
// \rfif.rdat2[7]~508_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\regs[24][7]~q )) # (!Instr_IF_19 & ((\regs[16][7]~q )))))

	.dataa(Instr_IF_18),
	.datab(\regs[24][7]~q ),
	.datac(\regs[16][7]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~508_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~508 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[7]~508 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N23
dffeas \regs[28][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][7] .is_wysiwyg = "true";
defparam \regs[28][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[7]~509 (
// Equation(s):
// \rfif.rdat2[7]~509_combout  = (\rfif.rdat2[7]~508_combout  & (((\regs[28][7]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[7]~508_combout  & (\regs[20][7]~q  & ((Instr_IF_18))))

	.dataa(\rfif.rdat2[7]~508_combout ),
	.datab(\regs[20][7]~q ),
	.datac(\regs[28][7]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~509_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~509 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[7]~509 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N13
dffeas \regs[24][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][6] .is_wysiwyg = "true";
defparam \regs[24][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N23
dffeas \regs[16][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][6] .is_wysiwyg = "true";
defparam \regs[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[6]~529 (
// Equation(s):
// \rfif.rdat2[6]~529_combout  = (Instr_IF_18 & ((\regs[20][6]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[16][6]~q  & !Instr_IF_19))))

	.dataa(\regs[20][6]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[16][6]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~529_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~529 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[6]~529 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \rfif.rdat2[6]~530 (
// Equation(s):
// \rfif.rdat2[6]~530_combout  = (\rfif.rdat2[6]~529_combout  & (((\regs[28][6]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[6]~529_combout  & (\regs[24][6]~q  & (Instr_IF_19)))

	.dataa(\regs[24][6]~q ),
	.datab(\rfif.rdat2[6]~529_combout ),
	.datac(Instr_IF_19),
	.datad(\regs[28][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~530_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~530 .lut_mask = 16'hEC2C;
defparam \rfif.rdat2[6]~530 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[6]~532 (
// Equation(s):
// \rfif.rdat2[6]~532_combout  = (Instr_IF_19 & ((\regs[27][6]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[19][6]~q  & !Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][6]~q ),
	.datac(\regs[19][6]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~532_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~532 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[6]~532 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \rfif.rdat2[6]~542 (
// Equation(s):
// \rfif.rdat2[6]~542_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][6]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][6]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][6]~q ),
	.datad(\regs[13][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~542_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~542 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[6]~542 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[6]~504 (
// Equation(s):
// \rfif.rdat1[6]~504_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][6]~q ))) # (!Instr_IF_24 & (\regs[16][6]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][6]~q ),
	.datac(\regs[24][6]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~504_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~504 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[6]~504 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[6]~512 (
// Equation(s):
// \rfif.rdat1[6]~512_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][6]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][6]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][6]~q ),
	.datad(\regs[4][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~512_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~512 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[6]~512 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[6]~514 (
// Equation(s):
// \rfif.rdat1[6]~514_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][6]~q )) # (!Instr_IF_21 & ((\regs[0][6]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][6]~q ),
	.datad(\regs[0][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~514_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~514 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[6]~514 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \regs[18][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][5] .is_wysiwyg = "true";
defparam \regs[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[5]~546 (
// Equation(s):
// \rfif.rdat2[5]~546_combout  = (Instr_IF_19 & (((\regs[26][5]~q ) # (Instr_IF_18)))) # (!Instr_IF_19 & (\regs[18][5]~q  & ((!Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[18][5]~q ),
	.datac(\regs[26][5]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~546_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~546 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[5]~546 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N27
dffeas \regs[17][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][5] .is_wysiwyg = "true";
defparam \regs[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[5]~548 (
// Equation(s):
// \rfif.rdat2[5]~548_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][5]~q ))) # (!Instr_IF_18 & (\regs[17][5]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][5]~q ),
	.datad(\regs[21][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~548_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~548 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[5]~548 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[5]~549 (
// Equation(s):
// \rfif.rdat2[5]~549_combout  = (\rfif.rdat2[5]~548_combout  & (((\regs[29][5]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[5]~548_combout  & (\regs[25][5]~q  & ((Instr_IF_19))))

	.dataa(\regs[25][5]~q ),
	.datab(\rfif.rdat2[5]~548_combout ),
	.datac(\regs[29][5]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~549_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~549 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[5]~549 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N13
dffeas \regs[20][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][5] .is_wysiwyg = "true";
defparam \regs[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[5]~553 (
// Equation(s):
// \rfif.rdat2[5]~553_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[23][5]~q )) # (!Instr_IF_18 & ((\regs[19][5]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[23][5]~q ),
	.datac(\regs[19][5]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~553_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~553 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[5]~553 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[5]~522 (
// Equation(s):
// \rfif.rdat1[5]~522_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[22][5]~q )) # (!Instr_IF_23 & ((\regs[18][5]~q )))))

	.dataa(Instr_IF_24),
	.datab(\regs[22][5]~q ),
	.datac(\regs[18][5]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~522_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~522 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[5]~522 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[5]~524 (
// Equation(s):
// \rfif.rdat1[5]~524_combout  = (Instr_IF_23 & (((\regs[20][5]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][5]~q  & ((!Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][5]~q ),
	.datac(\regs[20][5]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~524_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~524 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[5]~524 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N23
dffeas \regs[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][4] .is_wysiwyg = "true";
defparam \regs[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[4]~574 (
// Equation(s):
// \rfif.rdat2[4]~574_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[27][4]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[19][4]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][4]~q ),
	.datad(\regs[27][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~574_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~574 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[4]~574 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N16
cycloneive_lcell_comb \rfif.rdat2[4]~579 (
// Equation(s):
// \rfif.rdat2[4]~579_combout  = (Instr_IF_17 & (((Instr_IF_16) # (\regs[10][4]~q )))) # (!Instr_IF_17 & (\regs[8][4]~q  & (!Instr_IF_16)))

	.dataa(\regs[8][4]~q ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\regs[10][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~579_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~579 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[4]~579 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \rfif.rdat2[4]~580 (
// Equation(s):
// \rfif.rdat2[4]~580_combout  = (Instr_IF_16 & ((\rfif.rdat2[4]~579_combout  & ((\regs[11][4]~q ))) # (!\rfif.rdat2[4]~579_combout  & (\regs[9][4]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[4]~579_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][4]~q ),
	.datac(\regs[11][4]~q ),
	.datad(\rfif.rdat2[4]~579_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~580_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~580 .lut_mask = 16'hF588;
defparam \rfif.rdat2[4]~580 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N9
dffeas \regs[20][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][3] .is_wysiwyg = "true";
defparam \regs[20][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[3]~595 (
// Equation(s):
// \rfif.rdat2[3]~595_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[23][3]~q ))) # (!Instr_IF_18 & (\regs[19][3]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][3]~q ),
	.datad(\regs[23][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~595_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~595 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[3]~595 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[3]~598 (
// Equation(s):
// \rfif.rdat2[3]~598_combout  = (Instr_IF_16 & (((\regs[9][3]~q ) # (Instr_IF_17)))) # (!Instr_IF_16 & (\regs[8][3]~q  & ((!Instr_IF_17))))

	.dataa(\regs[8][3]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[9][3]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~598_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~598 .lut_mask = 16'hCCE2;
defparam \rfif.rdat2[3]~598 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N23
dffeas \regs[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][3] .is_wysiwyg = "true";
defparam \regs[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[3]~600 (
// Equation(s):
// \rfif.rdat2[3]~600_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][3]~q ))) # (!Instr_IF_17 & (\regs[4][3]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][3]~q ),
	.datad(\regs[6][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~600_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~600 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[3]~600 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[3]~601 (
// Equation(s):
// \rfif.rdat2[3]~601_combout  = (Instr_IF_16 & ((\rfif.rdat2[3]~600_combout  & (\regs[7][3]~q )) # (!\rfif.rdat2[3]~600_combout  & ((\regs[5][3]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[3]~600_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[3]~600_combout ),
	.datac(\regs[7][3]~q ),
	.datad(\regs[5][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~601_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~601 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[3]~601 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N31
dffeas \regs[0][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][3] .is_wysiwyg = "true";
defparam \regs[0][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[3]~602 (
// Equation(s):
// \rfif.rdat2[3]~602_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][3]~q ))) # (!Instr_IF_16 & (\regs[0][3]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][3]~q ),
	.datad(\regs[1][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~602_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~602 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[3]~602 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \rfif.rdat1[3]~562 (
// Equation(s):
// \rfif.rdat1[3]~562_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[22][3]~q )) # (!Instr_IF_23 & ((\regs[18][3]~q )))))

	.dataa(Instr_IF_24),
	.datab(\regs[22][3]~q ),
	.datac(\regs[18][3]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~562_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~562 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[3]~562 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[3]~564 (
// Equation(s):
// \rfif.rdat1[3]~564_combout  = (Instr_IF_23 & (((\regs[20][3]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][3]~q  & ((!Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][3]~q ),
	.datac(\regs[20][3]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~564_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~564 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[3]~564 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \regs[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][2] .is_wysiwyg = "true";
defparam \regs[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[2]~616 (
// Equation(s):
// \rfif.rdat2[2]~616_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[27][2]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[19][2]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][2]~q ),
	.datad(\regs[27][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~616_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~616 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[2]~616 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \rfif.rdat2[1]~630 (
// Equation(s):
// \rfif.rdat2[1]~630_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][1]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\regs[18][1]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[26][1]~q ),
	.datad(\regs[18][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~630_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~630 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[1]~630 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N31
dffeas \regs[16][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][1] .is_wysiwyg = "true";
defparam \regs[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N30
cycloneive_lcell_comb \rfif.rdat2[1]~634 (
// Equation(s):
// \rfif.rdat2[1]~634_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][1]~q ))) # (!Instr_IF_19 & (\regs[16][1]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][1]~q ),
	.datad(\regs[24][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~634_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~634 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[1]~634 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[1]~637 (
// Equation(s):
// \rfif.rdat2[1]~637_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[23][1]~q ))) # (!Instr_IF_18 & (\regs[19][1]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][1]~q ),
	.datad(\regs[23][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~637_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~637 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[1]~637 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[0]~653 (
// Equation(s):
// \rfif.rdat2[0]~653_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][0]~q ))) # (!Instr_IF_18 & (\regs[18][0]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][0]~q ),
	.datad(\regs[22][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~653_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~653 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[0]~653 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N27
dffeas \regs[16][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][0] .is_wysiwyg = "true";
defparam \regs[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[0]~655 (
// Equation(s):
// \rfif.rdat2[0]~655_combout  = (Instr_IF_18 & ((\regs[20][0]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[16][0]~q  & !Instr_IF_19))))

	.dataa(\regs[20][0]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[16][0]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~655_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~655 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[0]~655 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N31
dffeas \regs[19][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][0] .is_wysiwyg = "true";
defparam \regs[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[0]~658 (
// Equation(s):
// \rfif.rdat2[0]~658_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[27][0]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[19][0]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][0]~q ),
	.datad(\regs[27][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~658_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~658 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[0]~658 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \rfif.rdat2[0]~661 (
// Equation(s):
// \rfif.rdat2[0]~661_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][0]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & ((\regs[4][0]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[5][0]~q ),
	.datad(\regs[4][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~661_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~661 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[0]~661 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[0]~663 (
// Equation(s):
// \rfif.rdat2[0]~663_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[10][0]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[8][0]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[8][0]~q ),
	.datad(\regs[10][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~663_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~663 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[0]~663 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[0]~664 (
// Equation(s):
// \rfif.rdat2[0]~664_combout  = (Instr_IF_16 & ((\rfif.rdat2[0]~663_combout  & ((\regs[11][0]~q ))) # (!\rfif.rdat2[0]~663_combout  & (\regs[9][0]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[0]~663_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][0]~q ),
	.datac(\regs[11][0]~q ),
	.datad(\rfif.rdat2[0]~663_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~664_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~664 .lut_mask = 16'hF588;
defparam \rfif.rdat2[0]~664 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N12
cycloneive_lcell_comb \regs[20][31]~feeder (
// Equation(s):
// \regs[20][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[20][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \regs[1][31]~feeder (
// Equation(s):
// \regs[1][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[1][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N22
cycloneive_lcell_comb \regs[28][29]~feeder (
// Equation(s):
// \regs[28][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[28][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \regs[3][26]~feeder (
// Equation(s):
// \regs[3][26]~feeder_combout  = \input_b~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b4),
	.cin(gnd),
	.combout(\regs[3][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][26]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N6
cycloneive_lcell_comb \regs[28][25]~feeder (
// Equation(s):
// \regs[28][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b5),
	.cin(gnd),
	.combout(\regs[28][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \regs[3][24]~feeder (
// Equation(s):
// \regs[3][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[3][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \regs[28][24]~feeder (
// Equation(s):
// \regs[28][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[28][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \regs[28][23]~feeder (
// Equation(s):
// \regs[28][23]~feeder_combout  = \input_b~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][23]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \regs[24][21]~feeder (
// Equation(s):
// \regs[24][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b9),
	.cin(gnd),
	.combout(\regs[24][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \regs[1][19]~feeder (
// Equation(s):
// \regs[1][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b11),
	.cin(gnd),
	.combout(\regs[1][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \regs[2][19]~feeder (
// Equation(s):
// \regs[2][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \regs[3][16]~feeder (
// Equation(s):
// \regs[3][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b14),
	.cin(gnd),
	.combout(\regs[3][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \regs[7][12]~feeder (
// Equation(s):
// \regs[7][12]~feeder_combout  = \input_a~99_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a2),
	.cin(gnd),
	.combout(\regs[7][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[7][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N6
cycloneive_lcell_comb \regs[9][9]~feeder (
// Equation(s):
// \regs[9][9]~feeder_combout  = \input_a~108_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a5),
	.cin(gnd),
	.combout(\regs[9][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[31]~20 (
// Equation(s):
// rfifrdat2_31 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[31]~9_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[31]~19_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[31]~19_combout ),
	.datad(\rfif.rdat2[31]~9_combout ),
	.cin(gnd),
	.combout(rfifrdat2_31),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~20 .lut_mask = 16'hC840;
defparam \rfif.rdat2[31]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[31]~9 (
// Equation(s):
// rfifrdat1_31 = (Instr_IF_22 & ((\rfif.rdat1[31]~6_combout  & ((\rfif.rdat1[31]~8_combout ))) # (!\rfif.rdat1[31]~6_combout  & (\rfif.rdat1[31]~1_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[31]~6_combout ))))

	.dataa(\rfif.rdat1[31]~1_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[31]~8_combout ),
	.datad(\rfif.rdat1[31]~6_combout ),
	.cin(gnd),
	.combout(rfifrdat1_31),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~9 .lut_mask = 16'hF388;
defparam \rfif.rdat1[31]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[31]~19 (
// Equation(s):
// rfifrdat1_311 = (Instr_IF_24 & ((\rfif.rdat1[31]~16_combout  & ((\rfif.rdat1[31]~18_combout ))) # (!\rfif.rdat1[31]~16_combout  & (\rfif.rdat1[31]~11_combout )))) # (!Instr_IF_24 & (((\rfif.rdat1[31]~16_combout ))))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[31]~11_combout ),
	.datac(\rfif.rdat1[31]~16_combout ),
	.datad(\rfif.rdat1[31]~18_combout ),
	.cin(gnd),
	.combout(rfifrdat1_311),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~19 .lut_mask = 16'hF858;
defparam \rfif.rdat1[31]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \WideOr0~0 (
// Equation(s):
// WideOr0 = (Instr_IF_24) # ((Instr_IF_25) # ((Instr_IF_23) # (Instr_IF_22)))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_25),
	.datac(Instr_IF_23),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
// synopsys translate_off
defparam \WideOr0~0 .lut_mask = 16'hFFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \rfif.rdat1[30]~29 (
// Equation(s):
// rfifrdat1_30 = (Instr_IF_21 & ((\rfif.rdat1[30]~26_combout  & (\rfif.rdat1[30]~28_combout )) # (!\rfif.rdat1[30]~26_combout  & ((\rfif.rdat1[30]~21_combout ))))) # (!Instr_IF_21 & (((\rfif.rdat1[30]~26_combout ))))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[30]~28_combout ),
	.datac(\rfif.rdat1[30]~26_combout ),
	.datad(\rfif.rdat1[30]~21_combout ),
	.cin(gnd),
	.combout(rfifrdat1_30),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~29 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[30]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[30]~39 (
// Equation(s):
// rfifrdat1_301 = (\rfif.rdat1[30]~36_combout  & ((\rfif.rdat1[30]~38_combout ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[30]~36_combout  & (((\rfif.rdat1[30]~31_combout  & Instr_IF_23))))

	.dataa(\rfif.rdat1[30]~36_combout ),
	.datab(\rfif.rdat1[30]~38_combout ),
	.datac(\rfif.rdat1[30]~31_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(rfifrdat1_301),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~39 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[30]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \rfif.rdat2[30]~41 (
// Equation(s):
// rfifrdat2_30 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[30]~30_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[30]~40_combout ))))

	.dataa(\rfif.rdat2[30]~40_combout ),
	.datab(Instr_IF_20),
	.datac(\WideOr1~combout ),
	.datad(\rfif.rdat2[30]~30_combout ),
	.cin(gnd),
	.combout(rfifrdat2_30),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~41 .lut_mask = 16'hE020;
defparam \rfif.rdat2[30]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \rfif.rdat1[29]~49 (
// Equation(s):
// rfifrdat1_29 = (Instr_IF_22 & ((\rfif.rdat1[29]~46_combout  & ((\rfif.rdat1[29]~48_combout ))) # (!\rfif.rdat1[29]~46_combout  & (\rfif.rdat1[29]~41_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[29]~46_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[29]~41_combout ),
	.datac(\rfif.rdat1[29]~46_combout ),
	.datad(\rfif.rdat1[29]~48_combout ),
	.cin(gnd),
	.combout(rfifrdat1_29),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~49 .lut_mask = 16'hF858;
defparam \rfif.rdat1[29]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[29]~59 (
// Equation(s):
// rfifrdat1_291 = (\rfif.rdat1[29]~56_combout  & ((\rfif.rdat1[29]~58_combout ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[29]~56_combout  & (((Instr_IF_24 & \rfif.rdat1[29]~51_combout ))))

	.dataa(\rfif.rdat1[29]~58_combout ),
	.datab(\rfif.rdat1[29]~56_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[29]~51_combout ),
	.cin(gnd),
	.combout(rfifrdat1_291),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~59 .lut_mask = 16'hBC8C;
defparam \rfif.rdat1[29]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \rfif.rdat2[29]~62 (
// Equation(s):
// rfifrdat2_29 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[29]~51_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[29]~61_combout ))))

	.dataa(\rfif.rdat2[29]~61_combout ),
	.datab(\WideOr1~combout ),
	.datac(Instr_IF_20),
	.datad(\rfif.rdat2[29]~51_combout ),
	.cin(gnd),
	.combout(rfifrdat2_29),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~62 .lut_mask = 16'hC808;
defparam \rfif.rdat2[29]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \rfif.rdat1[28]~69 (
// Equation(s):
// rfifrdat1_28 = (Instr_IF_21 & ((\rfif.rdat1[28]~66_combout  & (\rfif.rdat1[28]~68_combout )) # (!\rfif.rdat1[28]~66_combout  & ((\rfif.rdat1[28]~61_combout ))))) # (!Instr_IF_21 & (\rfif.rdat1[28]~66_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[28]~66_combout ),
	.datac(\rfif.rdat1[28]~68_combout ),
	.datad(\rfif.rdat1[28]~61_combout ),
	.cin(gnd),
	.combout(rfifrdat1_28),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~69 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[28]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \rfif.rdat1[28]~79 (
// Equation(s):
// rfifrdat1_281 = (Instr_IF_23 & ((\rfif.rdat1[28]~76_combout  & (\rfif.rdat1[28]~78_combout )) # (!\rfif.rdat1[28]~76_combout  & ((\rfif.rdat1[28]~71_combout ))))) # (!Instr_IF_23 & (((\rfif.rdat1[28]~76_combout ))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[28]~78_combout ),
	.datac(\rfif.rdat1[28]~76_combout ),
	.datad(\rfif.rdat1[28]~71_combout ),
	.cin(gnd),
	.combout(rfifrdat1_281),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~79 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[28]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[28]~83 (
// Equation(s):
// rfifrdat2_28 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[28]~72_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[28]~82_combout ))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[28]~82_combout ),
	.datad(\rfif.rdat2[28]~72_combout ),
	.cin(gnd),
	.combout(rfifrdat2_28),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~83 .lut_mask = 16'hA820;
defparam \rfif.rdat2[28]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[27]~89 (
// Equation(s):
// rfifrdat1_27 = (Instr_IF_22 & ((\rfif.rdat1[27]~86_combout  & (\rfif.rdat1[27]~88_combout )) # (!\rfif.rdat1[27]~86_combout  & ((\rfif.rdat1[27]~81_combout ))))) # (!Instr_IF_22 & (((\rfif.rdat1[27]~86_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[27]~88_combout ),
	.datac(\rfif.rdat1[27]~81_combout ),
	.datad(\rfif.rdat1[27]~86_combout ),
	.cin(gnd),
	.combout(rfifrdat1_27),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~89 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[27]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \rfif.rdat1[27]~99 (
// Equation(s):
// rfifrdat1_271 = (\rfif.rdat1[27]~96_combout  & ((\rfif.rdat1[27]~98_combout ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[27]~96_combout  & (((Instr_IF_24 & \rfif.rdat1[27]~91_combout ))))

	.dataa(\rfif.rdat1[27]~96_combout ),
	.datab(\rfif.rdat1[27]~98_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[27]~91_combout ),
	.cin(gnd),
	.combout(rfifrdat1_271),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~99 .lut_mask = 16'hDA8A;
defparam \rfif.rdat1[27]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \rfif.rdat2[27]~104 (
// Equation(s):
// rfifrdat2_27 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[27]~93_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[27]~103_combout ))))

	.dataa(\rfif.rdat2[27]~103_combout ),
	.datab(\WideOr1~combout ),
	.datac(Instr_IF_20),
	.datad(\rfif.rdat2[27]~93_combout ),
	.cin(gnd),
	.combout(rfifrdat2_27),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~104 .lut_mask = 16'hC808;
defparam \rfif.rdat2[27]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \rfif.rdat1[26]~109 (
// Equation(s):
// rfifrdat1_26 = (Instr_IF_21 & ((\rfif.rdat1[26]~106_combout  & (\rfif.rdat1[26]~108_combout )) # (!\rfif.rdat1[26]~106_combout  & ((\rfif.rdat1[26]~101_combout ))))) # (!Instr_IF_21 & (((\rfif.rdat1[26]~106_combout ))))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[26]~108_combout ),
	.datac(\rfif.rdat1[26]~101_combout ),
	.datad(\rfif.rdat1[26]~106_combout ),
	.cin(gnd),
	.combout(rfifrdat1_26),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~109 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[26]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \rfif.rdat1[26]~119 (
// Equation(s):
// rfifrdat1_261 = (Instr_IF_23 & ((\rfif.rdat1[26]~116_combout  & ((\rfif.rdat1[26]~118_combout ))) # (!\rfif.rdat1[26]~116_combout  & (\rfif.rdat1[26]~111_combout )))) # (!Instr_IF_23 & (((\rfif.rdat1[26]~116_combout ))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[26]~111_combout ),
	.datac(\rfif.rdat1[26]~118_combout ),
	.datad(\rfif.rdat1[26]~116_combout ),
	.cin(gnd),
	.combout(rfifrdat1_261),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~119 .lut_mask = 16'hF588;
defparam \rfif.rdat1[26]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \rfif.rdat2[26]~125 (
// Equation(s):
// rfifrdat2_26 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[26]~114_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[26]~124_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[26]~124_combout ),
	.datad(\rfif.rdat2[26]~114_combout ),
	.cin(gnd),
	.combout(rfifrdat2_26),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~125 .lut_mask = 16'hC840;
defparam \rfif.rdat2[26]~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \rfif.rdat1[25]~129 (
// Equation(s):
// rfifrdat1_25 = (Instr_IF_22 & ((\rfif.rdat1[25]~126_combout  & (\rfif.rdat1[25]~128_combout )) # (!\rfif.rdat1[25]~126_combout  & ((\rfif.rdat1[25]~121_combout ))))) # (!Instr_IF_22 & (((\rfif.rdat1[25]~126_combout ))))

	.dataa(\rfif.rdat1[25]~128_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[25]~121_combout ),
	.datad(\rfif.rdat1[25]~126_combout ),
	.cin(gnd),
	.combout(rfifrdat1_25),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~129 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[25]~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \rfif.rdat1[25]~139 (
// Equation(s):
// rfifrdat1_251 = (\rfif.rdat1[25]~136_combout  & (((\rfif.rdat1[25]~138_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[25]~136_combout  & (\rfif.rdat1[25]~131_combout  & (Instr_IF_24)))

	.dataa(\rfif.rdat1[25]~136_combout ),
	.datab(\rfif.rdat1[25]~131_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[25]~138_combout ),
	.cin(gnd),
	.combout(rfifrdat1_251),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~139 .lut_mask = 16'hEA4A;
defparam \rfif.rdat1[25]~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[25]~146 (
// Equation(s):
// rfifrdat2_25 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[25]~135_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[25]~145_combout ))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[25]~145_combout ),
	.datad(\rfif.rdat2[25]~135_combout ),
	.cin(gnd),
	.combout(rfifrdat2_25),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~146 .lut_mask = 16'hA820;
defparam \rfif.rdat2[25]~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \rfif.rdat1[24]~149 (
// Equation(s):
// rfifrdat1_24 = (\rfif.rdat1[24]~146_combout  & (((\rfif.rdat1[24]~148_combout ) # (!Instr_IF_21)))) # (!\rfif.rdat1[24]~146_combout  & (\rfif.rdat1[24]~141_combout  & (Instr_IF_21)))

	.dataa(\rfif.rdat1[24]~141_combout ),
	.datab(\rfif.rdat1[24]~146_combout ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[24]~148_combout ),
	.cin(gnd),
	.combout(rfifrdat1_24),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~149 .lut_mask = 16'hEC2C;
defparam \rfif.rdat1[24]~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \rfif.rdat1[24]~159 (
// Equation(s):
// rfifrdat1_241 = (Instr_IF_23 & ((\rfif.rdat1[24]~156_combout  & (\rfif.rdat1[24]~158_combout )) # (!\rfif.rdat1[24]~156_combout  & ((\rfif.rdat1[24]~151_combout ))))) # (!Instr_IF_23 & (((\rfif.rdat1[24]~156_combout ))))

	.dataa(\rfif.rdat1[24]~158_combout ),
	.datab(\rfif.rdat1[24]~151_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[24]~156_combout ),
	.cin(gnd),
	.combout(rfifrdat1_241),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~159 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[24]~159 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \rfif.rdat2[24]~167 (
// Equation(s):
// rfifrdat2_24 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[24]~156_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[24]~166_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[24]~156_combout ),
	.datad(\rfif.rdat2[24]~166_combout ),
	.cin(gnd),
	.combout(rfifrdat2_24),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~167 .lut_mask = 16'hA280;
defparam \rfif.rdat2[24]~167 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[23]~169 (
// Equation(s):
// rfifrdat1_23 = (Instr_IF_22 & ((\rfif.rdat1[23]~166_combout  & ((\rfif.rdat1[23]~168_combout ))) # (!\rfif.rdat1[23]~166_combout  & (\rfif.rdat1[23]~161_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[23]~166_combout ))))

	.dataa(\rfif.rdat1[23]~161_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[23]~168_combout ),
	.datad(\rfif.rdat1[23]~166_combout ),
	.cin(gnd),
	.combout(rfifrdat1_23),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~169 .lut_mask = 16'hF388;
defparam \rfif.rdat1[23]~169 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[23]~179 (
// Equation(s):
// rfifrdat1_231 = (Instr_IF_24 & ((\rfif.rdat1[23]~176_combout  & (\rfif.rdat1[23]~178_combout )) # (!\rfif.rdat1[23]~176_combout  & ((\rfif.rdat1[23]~171_combout ))))) # (!Instr_IF_24 & (\rfif.rdat1[23]~176_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[23]~176_combout ),
	.datac(\rfif.rdat1[23]~178_combout ),
	.datad(\rfif.rdat1[23]~171_combout ),
	.cin(gnd),
	.combout(rfifrdat1_231),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~179 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[23]~179 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \rfif.rdat2[23]~188 (
// Equation(s):
// rfifrdat2_23 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[23]~177_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[23]~187_combout ))))

	.dataa(\rfif.rdat2[23]~187_combout ),
	.datab(Instr_IF_20),
	.datac(\WideOr1~combout ),
	.datad(\rfif.rdat2[23]~177_combout ),
	.cin(gnd),
	.combout(rfifrdat2_23),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~188 .lut_mask = 16'hE020;
defparam \rfif.rdat2[23]~188 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \rfif.rdat1[22]~189 (
// Equation(s):
// rfifrdat1_22 = (Instr_IF_21 & ((\rfif.rdat1[22]~186_combout  & ((\rfif.rdat1[22]~188_combout ))) # (!\rfif.rdat1[22]~186_combout  & (\rfif.rdat1[22]~181_combout )))) # (!Instr_IF_21 & (\rfif.rdat1[22]~186_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[22]~186_combout ),
	.datac(\rfif.rdat1[22]~181_combout ),
	.datad(\rfif.rdat1[22]~188_combout ),
	.cin(gnd),
	.combout(rfifrdat1_22),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~189 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[22]~189 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \rfif.rdat1[22]~199 (
// Equation(s):
// rfifrdat1_221 = (\rfif.rdat1[22]~196_combout  & ((\rfif.rdat1[22]~198_combout ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[22]~196_combout  & (((\rfif.rdat1[22]~191_combout  & Instr_IF_23))))

	.dataa(\rfif.rdat1[22]~198_combout ),
	.datab(\rfif.rdat1[22]~196_combout ),
	.datac(\rfif.rdat1[22]~191_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(rfifrdat1_221),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~199 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[22]~199 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \rfif.rdat2[22]~209 (
// Equation(s):
// rfifrdat2_22 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[22]~198_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[22]~208_combout )))))

	.dataa(\rfif.rdat2[22]~198_combout ),
	.datab(\rfif.rdat2[22]~208_combout ),
	.datac(\WideOr1~combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_22),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~209 .lut_mask = 16'hA0C0;
defparam \rfif.rdat2[22]~209 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \rfif.rdat1[21]~209 (
// Equation(s):
// rfifrdat1_21 = (\rfif.rdat1[21]~206_combout  & ((\rfif.rdat1[21]~208_combout ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[21]~206_combout  & (((Instr_IF_22 & \rfif.rdat1[21]~201_combout ))))

	.dataa(\rfif.rdat1[21]~206_combout ),
	.datab(\rfif.rdat1[21]~208_combout ),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[21]~201_combout ),
	.cin(gnd),
	.combout(rfifrdat1_21),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~209 .lut_mask = 16'hDA8A;
defparam \rfif.rdat1[21]~209 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \rfif.rdat1[21]~219 (
// Equation(s):
// rfifrdat1_211 = (\rfif.rdat1[21]~216_combout  & (((\rfif.rdat1[21]~218_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[21]~216_combout  & (\rfif.rdat1[21]~211_combout  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[21]~216_combout ),
	.datab(\rfif.rdat1[21]~211_combout ),
	.datac(\rfif.rdat1[21]~218_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_211),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~219 .lut_mask = 16'hE4AA;
defparam \rfif.rdat1[21]~219 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \rfif.rdat2[21]~230 (
// Equation(s):
// rfifrdat2_21 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[21]~219_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[21]~229_combout ))))

	.dataa(\rfif.rdat2[21]~229_combout ),
	.datab(\WideOr1~combout ),
	.datac(Instr_IF_20),
	.datad(\rfif.rdat2[21]~219_combout ),
	.cin(gnd),
	.combout(rfifrdat2_21),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~230 .lut_mask = 16'hC808;
defparam \rfif.rdat2[21]~230 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[20]~229 (
// Equation(s):
// rfifrdat1_20 = (Instr_IF_21 & ((\rfif.rdat1[20]~226_combout  & (\rfif.rdat1[20]~228_combout )) # (!\rfif.rdat1[20]~226_combout  & ((\rfif.rdat1[20]~221_combout ))))) # (!Instr_IF_21 & (((\rfif.rdat1[20]~226_combout ))))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[20]~228_combout ),
	.datac(\rfif.rdat1[20]~221_combout ),
	.datad(\rfif.rdat1[20]~226_combout ),
	.cin(gnd),
	.combout(rfifrdat1_20),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~229 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[20]~229 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[20]~239 (
// Equation(s):
// rfifrdat1_201 = (\rfif.rdat1[20]~236_combout  & (((\rfif.rdat1[20]~238_combout )) # (!Instr_IF_23))) # (!\rfif.rdat1[20]~236_combout  & (Instr_IF_23 & ((\rfif.rdat1[20]~231_combout ))))

	.dataa(\rfif.rdat1[20]~236_combout ),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[20]~238_combout ),
	.datad(\rfif.rdat1[20]~231_combout ),
	.cin(gnd),
	.combout(rfifrdat1_201),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~239 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[20]~239 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \rfif.rdat2[20]~251 (
// Equation(s):
// rfifrdat2_20 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[20]~240_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[20]~250_combout )))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[20]~240_combout ),
	.datad(\rfif.rdat2[20]~250_combout ),
	.cin(gnd),
	.combout(rfifrdat2_20),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~251 .lut_mask = 16'hC480;
defparam \rfif.rdat2[20]~251 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[19]~249 (
// Equation(s):
// rfifrdat1_19 = (Instr_IF_22 & ((\rfif.rdat1[19]~246_combout  & ((\rfif.rdat1[19]~248_combout ))) # (!\rfif.rdat1[19]~246_combout  & (\rfif.rdat1[19]~241_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[19]~246_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[19]~241_combout ),
	.datac(\rfif.rdat1[19]~248_combout ),
	.datad(\rfif.rdat1[19]~246_combout ),
	.cin(gnd),
	.combout(rfifrdat1_19),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~249 .lut_mask = 16'hF588;
defparam \rfif.rdat1[19]~249 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \rfif.rdat1[19]~259 (
// Equation(s):
// rfifrdat1_191 = (\rfif.rdat1[19]~256_combout  & (((\rfif.rdat1[19]~258_combout )) # (!Instr_IF_24))) # (!\rfif.rdat1[19]~256_combout  & (Instr_IF_24 & (\rfif.rdat1[19]~251_combout )))

	.dataa(\rfif.rdat1[19]~256_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[19]~251_combout ),
	.datad(\rfif.rdat1[19]~258_combout ),
	.cin(gnd),
	.combout(rfifrdat1_191),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~259 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[19]~259 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \rfif.rdat2[19]~272 (
// Equation(s):
// rfifrdat2_19 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[19]~261_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[19]~271_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[19]~271_combout ),
	.datad(\rfif.rdat2[19]~261_combout ),
	.cin(gnd),
	.combout(rfifrdat2_19),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~272 .lut_mask = 16'hC840;
defparam \rfif.rdat2[19]~272 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[18]~269 (
// Equation(s):
// rfifrdat1_18 = (Instr_IF_21 & ((\rfif.rdat1[18]~266_combout  & ((\rfif.rdat1[18]~268_combout ))) # (!\rfif.rdat1[18]~266_combout  & (\rfif.rdat1[18]~261_combout )))) # (!Instr_IF_21 & (((\rfif.rdat1[18]~266_combout ))))

	.dataa(\rfif.rdat1[18]~261_combout ),
	.datab(\rfif.rdat1[18]~268_combout ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[18]~266_combout ),
	.cin(gnd),
	.combout(rfifrdat1_18),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~269 .lut_mask = 16'hCFA0;
defparam \rfif.rdat1[18]~269 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \rfif.rdat1[18]~279 (
// Equation(s):
// rfifrdat1_181 = (Instr_IF_23 & ((\rfif.rdat1[18]~276_combout  & (\rfif.rdat1[18]~278_combout )) # (!\rfif.rdat1[18]~276_combout  & ((\rfif.rdat1[18]~271_combout ))))) # (!Instr_IF_23 & (((\rfif.rdat1[18]~276_combout ))))

	.dataa(\rfif.rdat1[18]~278_combout ),
	.datab(\rfif.rdat1[18]~271_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[18]~276_combout ),
	.cin(gnd),
	.combout(rfifrdat1_181),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~279 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[18]~279 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \rfif.rdat2[18]~293 (
// Equation(s):
// rfifrdat2_18 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[18]~282_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[18]~292_combout )))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[18]~282_combout ),
	.datad(\rfif.rdat2[18]~292_combout ),
	.cin(gnd),
	.combout(rfifrdat2_18),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~293 .lut_mask = 16'hC480;
defparam \rfif.rdat2[18]~293 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \rfif.rdat1[17]~289 (
// Equation(s):
// rfifrdat1_17 = (Instr_IF_22 & ((\rfif.rdat1[17]~286_combout  & ((\rfif.rdat1[17]~288_combout ))) # (!\rfif.rdat1[17]~286_combout  & (\rfif.rdat1[17]~281_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[17]~286_combout ))))

	.dataa(\rfif.rdat1[17]~281_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[17]~286_combout ),
	.datad(\rfif.rdat1[17]~288_combout ),
	.cin(gnd),
	.combout(rfifrdat1_17),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~289 .lut_mask = 16'hF838;
defparam \rfif.rdat1[17]~289 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[17]~299 (
// Equation(s):
// rfifrdat1_171 = (Instr_IF_24 & ((\rfif.rdat1[17]~296_combout  & (\rfif.rdat1[17]~298_combout )) # (!\rfif.rdat1[17]~296_combout  & ((\rfif.rdat1[17]~291_combout ))))) # (!Instr_IF_24 & (((\rfif.rdat1[17]~296_combout ))))

	.dataa(\rfif.rdat1[17]~298_combout ),
	.datab(\rfif.rdat1[17]~291_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[17]~296_combout ),
	.cin(gnd),
	.combout(rfifrdat1_171),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~299 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[17]~299 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \rfif.rdat2[17]~314 (
// Equation(s):
// rfifrdat2_17 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[17]~303_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[17]~313_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[17]~303_combout ),
	.datad(\rfif.rdat2[17]~313_combout ),
	.cin(gnd),
	.combout(rfifrdat2_17),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~314 .lut_mask = 16'hA280;
defparam \rfif.rdat2[17]~314 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[16]~309 (
// Equation(s):
// rfifrdat1_16 = (Instr_IF_21 & ((\rfif.rdat1[16]~306_combout  & (\rfif.rdat1[16]~308_combout )) # (!\rfif.rdat1[16]~306_combout  & ((\rfif.rdat1[16]~301_combout ))))) # (!Instr_IF_21 & (((\rfif.rdat1[16]~306_combout ))))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[16]~308_combout ),
	.datac(\rfif.rdat1[16]~306_combout ),
	.datad(\rfif.rdat1[16]~301_combout ),
	.cin(gnd),
	.combout(rfifrdat1_16),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~309 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[16]~309 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[16]~319 (
// Equation(s):
// rfifrdat1_161 = (\rfif.rdat1[16]~316_combout  & (((\rfif.rdat1[16]~318_combout ) # (!Instr_IF_23)))) # (!\rfif.rdat1[16]~316_combout  & (\rfif.rdat1[16]~311_combout  & (Instr_IF_23)))

	.dataa(\rfif.rdat1[16]~316_combout ),
	.datab(\rfif.rdat1[16]~311_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[16]~318_combout ),
	.cin(gnd),
	.combout(rfifrdat1_161),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~319 .lut_mask = 16'hEA4A;
defparam \rfif.rdat1[16]~319 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \rfif.rdat2[16]~335 (
// Equation(s):
// rfifrdat2_16 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[16]~324_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[16]~334_combout ))))

	.dataa(\rfif.rdat2[16]~334_combout ),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[16]~324_combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_16),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~335 .lut_mask = 16'hC088;
defparam \rfif.rdat2[16]~335 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \rfif.rdat1[15]~329 (
// Equation(s):
// rfifrdat1_15 = (Instr_IF_22 & ((\rfif.rdat1[15]~326_combout  & ((\rfif.rdat1[15]~328_combout ))) # (!\rfif.rdat1[15]~326_combout  & (\rfif.rdat1[15]~321_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[15]~326_combout ))))

	.dataa(\rfif.rdat1[15]~321_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[15]~326_combout ),
	.datad(\rfif.rdat1[15]~328_combout ),
	.cin(gnd),
	.combout(rfifrdat1_15),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~329 .lut_mask = 16'hF838;
defparam \rfif.rdat1[15]~329 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[15]~339 (
// Equation(s):
// rfifrdat1_151 = (\rfif.rdat1[15]~336_combout  & (((\rfif.rdat1[15]~338_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[15]~336_combout  & (\rfif.rdat1[15]~331_combout  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[15]~331_combout ),
	.datab(\rfif.rdat1[15]~336_combout ),
	.datac(\rfif.rdat1[15]~338_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_151),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~339 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[15]~339 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[15]~356 (
// Equation(s):
// rfifrdat2_15 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[15]~345_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[15]~355_combout ))))

	.dataa(\rfif.rdat2[15]~355_combout ),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[15]~345_combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_15),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~356 .lut_mask = 16'hC088;
defparam \rfif.rdat2[15]~356 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \rfif.rdat1[14]~349 (
// Equation(s):
// rfifrdat1_14 = (Instr_IF_21 & ((\rfif.rdat1[14]~346_combout  & ((\rfif.rdat1[14]~348_combout ))) # (!\rfif.rdat1[14]~346_combout  & (\rfif.rdat1[14]~341_combout )))) # (!Instr_IF_21 & (((\rfif.rdat1[14]~346_combout ))))

	.dataa(\rfif.rdat1[14]~341_combout ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[14]~348_combout ),
	.datad(\rfif.rdat1[14]~346_combout ),
	.cin(gnd),
	.combout(rfifrdat1_14),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~349 .lut_mask = 16'hF388;
defparam \rfif.rdat1[14]~349 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[14]~359 (
// Equation(s):
// rfifrdat1_141 = (Instr_IF_23 & ((\rfif.rdat1[14]~356_combout  & (\rfif.rdat1[14]~358_combout )) # (!\rfif.rdat1[14]~356_combout  & ((\rfif.rdat1[14]~351_combout ))))) # (!Instr_IF_23 & (((\rfif.rdat1[14]~356_combout ))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[14]~358_combout ),
	.datac(\rfif.rdat1[14]~351_combout ),
	.datad(\rfif.rdat1[14]~356_combout ),
	.cin(gnd),
	.combout(rfifrdat1_141),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~359 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[14]~359 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N6
cycloneive_lcell_comb \rfif.rdat2[14]~377 (
// Equation(s):
// rfifrdat2_14 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[14]~366_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[14]~376_combout )))))

	.dataa(\rfif.rdat2[14]~366_combout ),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[14]~376_combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_14),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~377 .lut_mask = 16'h88C0;
defparam \rfif.rdat2[14]~377 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[13]~398 (
// Equation(s):
// rfifrdat2_13 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[13]~387_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[13]~397_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[13]~387_combout ),
	.datad(\rfif.rdat2[13]~397_combout ),
	.cin(gnd),
	.combout(rfifrdat2_13),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~398 .lut_mask = 16'hA280;
defparam \rfif.rdat2[13]~398 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[13]~369 (
// Equation(s):
// rfifrdat1_13 = (\rfif.rdat1[13]~366_combout  & (((\rfif.rdat1[13]~368_combout )) # (!Instr_IF_21))) # (!\rfif.rdat1[13]~366_combout  & (Instr_IF_21 & (\rfif.rdat1[13]~361_combout )))

	.dataa(\rfif.rdat1[13]~366_combout ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[13]~361_combout ),
	.datad(\rfif.rdat1[13]~368_combout ),
	.cin(gnd),
	.combout(rfifrdat1_13),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~369 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[13]~369 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[13]~379 (
// Equation(s):
// rfifrdat1_131 = (Instr_IF_23 & ((\rfif.rdat1[13]~376_combout  & ((\rfif.rdat1[13]~378_combout ))) # (!\rfif.rdat1[13]~376_combout  & (\rfif.rdat1[13]~371_combout )))) # (!Instr_IF_23 & (((\rfif.rdat1[13]~376_combout ))))

	.dataa(\rfif.rdat1[13]~371_combout ),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[13]~378_combout ),
	.datad(\rfif.rdat1[13]~376_combout ),
	.cin(gnd),
	.combout(rfifrdat1_131),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~379 .lut_mask = 16'hF388;
defparam \rfif.rdat1[13]~379 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[12]~419 (
// Equation(s):
// rfifrdat2_12 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[12]~408_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[12]~418_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[12]~408_combout ),
	.datad(\rfif.rdat2[12]~418_combout ),
	.cin(gnd),
	.combout(rfifrdat2_12),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~419 .lut_mask = 16'hA280;
defparam \rfif.rdat2[12]~419 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N10
cycloneive_lcell_comb \rfif.rdat1[12]~389 (
// Equation(s):
// rfifrdat1_12 = (Instr_IF_22 & ((\rfif.rdat1[12]~386_combout  & (\rfif.rdat1[12]~388_combout )) # (!\rfif.rdat1[12]~386_combout  & ((\rfif.rdat1[12]~381_combout ))))) # (!Instr_IF_22 & (\rfif.rdat1[12]~386_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[12]~386_combout ),
	.datac(\rfif.rdat1[12]~388_combout ),
	.datad(\rfif.rdat1[12]~381_combout ),
	.cin(gnd),
	.combout(rfifrdat1_12),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~389 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[12]~389 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N22
cycloneive_lcell_comb \rfif.rdat1[12]~399 (
// Equation(s):
// rfifrdat1_121 = (\rfif.rdat1[12]~396_combout  & (((\rfif.rdat1[12]~398_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[12]~396_combout  & (\rfif.rdat1[12]~391_combout  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[12]~391_combout ),
	.datab(\rfif.rdat1[12]~396_combout ),
	.datac(\rfif.rdat1[12]~398_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_121),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~399 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[12]~399 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[11]~440 (
// Equation(s):
// rfifrdat2_11 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[11]~429_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[11]~439_combout ))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[11]~439_combout ),
	.datad(\rfif.rdat2[11]~429_combout ),
	.cin(gnd),
	.combout(rfifrdat2_11),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~440 .lut_mask = 16'hA820;
defparam \rfif.rdat2[11]~440 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \rfif.rdat1[11]~409 (
// Equation(s):
// rfifrdat1_11 = (\rfif.rdat1[11]~406_combout  & ((\rfif.rdat1[11]~408_combout ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[11]~406_combout  & (((\rfif.rdat1[11]~401_combout  & Instr_IF_21))))

	.dataa(\rfif.rdat1[11]~408_combout ),
	.datab(\rfif.rdat1[11]~401_combout ),
	.datac(\rfif.rdat1[11]~406_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(rfifrdat1_11),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~409 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[11]~409 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \rfif.rdat1[11]~419 (
// Equation(s):
// rfifrdat1_111 = (\rfif.rdat1[11]~416_combout  & ((\rfif.rdat1[11]~418_combout ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[11]~416_combout  & (((\rfif.rdat1[11]~411_combout  & Instr_IF_23))))

	.dataa(\rfif.rdat1[11]~418_combout ),
	.datab(\rfif.rdat1[11]~416_combout ),
	.datac(\rfif.rdat1[11]~411_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(rfifrdat1_111),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~419 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[11]~419 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \rfif.rdat2[10]~461 (
// Equation(s):
// rfifrdat2_10 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[10]~450_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[10]~460_combout ))))

	.dataa(\rfif.rdat2[10]~460_combout ),
	.datab(Instr_IF_20),
	.datac(\WideOr1~combout ),
	.datad(\rfif.rdat2[10]~450_combout ),
	.cin(gnd),
	.combout(rfifrdat2_10),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~461 .lut_mask = 16'hE020;
defparam \rfif.rdat2[10]~461 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[10]~429 (
// Equation(s):
// rfifrdat1_10 = (Instr_IF_22 & ((\rfif.rdat1[10]~426_combout  & (\rfif.rdat1[10]~428_combout )) # (!\rfif.rdat1[10]~426_combout  & ((\rfif.rdat1[10]~421_combout ))))) # (!Instr_IF_22 & (((\rfif.rdat1[10]~426_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[10]~428_combout ),
	.datac(\rfif.rdat1[10]~421_combout ),
	.datad(\rfif.rdat1[10]~426_combout ),
	.cin(gnd),
	.combout(rfifrdat1_10),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~429 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[10]~429 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[10]~439 (
// Equation(s):
// rfifrdat1_101 = (\rfif.rdat1[10]~436_combout  & ((\rfif.rdat1[10]~438_combout ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[10]~436_combout  & (((\rfif.rdat1[10]~431_combout  & Instr_IF_24))))

	.dataa(\rfif.rdat1[10]~438_combout ),
	.datab(\rfif.rdat1[10]~436_combout ),
	.datac(\rfif.rdat1[10]~431_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_101),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~439 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[10]~439 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[9]~482 (
// Equation(s):
// rfifrdat2_9 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[9]~471_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[9]~481_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(\rfif.rdat2[9]~471_combout ),
	.datac(\rfif.rdat2[9]~481_combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_9),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~482 .lut_mask = 16'h88A0;
defparam \rfif.rdat2[9]~482 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[9]~449 (
// Equation(s):
// rfifrdat1_9 = (Instr_IF_21 & ((\rfif.rdat1[9]~446_combout  & ((\rfif.rdat1[9]~448_combout ))) # (!\rfif.rdat1[9]~446_combout  & (\rfif.rdat1[9]~441_combout )))) # (!Instr_IF_21 & (((\rfif.rdat1[9]~446_combout ))))

	.dataa(\rfif.rdat1[9]~441_combout ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[9]~448_combout ),
	.datad(\rfif.rdat1[9]~446_combout ),
	.cin(gnd),
	.combout(rfifrdat1_9),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~449 .lut_mask = 16'hF388;
defparam \rfif.rdat1[9]~449 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \rfif.rdat1[9]~459 (
// Equation(s):
// rfifrdat1_91 = (Instr_IF_23 & ((\rfif.rdat1[9]~456_combout  & (\rfif.rdat1[9]~458_combout )) # (!\rfif.rdat1[9]~456_combout  & ((\rfif.rdat1[9]~451_combout ))))) # (!Instr_IF_23 & (\rfif.rdat1[9]~456_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[9]~456_combout ),
	.datac(\rfif.rdat1[9]~458_combout ),
	.datad(\rfif.rdat1[9]~451_combout ),
	.cin(gnd),
	.combout(rfifrdat1_91),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~459 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[9]~459 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \rfif.rdat2[8]~503 (
// Equation(s):
// rfifrdat2_8 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[8]~492_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[8]~502_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(Instr_IF_20),
	.datac(\rfif.rdat2[8]~492_combout ),
	.datad(\rfif.rdat2[8]~502_combout ),
	.cin(gnd),
	.combout(rfifrdat2_8),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~503 .lut_mask = 16'hA280;
defparam \rfif.rdat2[8]~503 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \rfif.rdat1[8]~469 (
// Equation(s):
// rfifrdat1_8 = (Instr_IF_22 & ((\rfif.rdat1[8]~466_combout  & ((\rfif.rdat1[8]~468_combout ))) # (!\rfif.rdat1[8]~466_combout  & (\rfif.rdat1[8]~461_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[8]~466_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[8]~461_combout ),
	.datac(\rfif.rdat1[8]~466_combout ),
	.datad(\rfif.rdat1[8]~468_combout ),
	.cin(gnd),
	.combout(rfifrdat1_8),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~469 .lut_mask = 16'hF858;
defparam \rfif.rdat1[8]~469 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[8]~479 (
// Equation(s):
// rfifrdat1_81 = (\rfif.rdat1[8]~476_combout  & (((\rfif.rdat1[8]~478_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[8]~476_combout  & (\rfif.rdat1[8]~471_combout  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[8]~471_combout ),
	.datab(\rfif.rdat1[8]~478_combout ),
	.datac(\rfif.rdat1[8]~476_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_81),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~479 .lut_mask = 16'hCAF0;
defparam \rfif.rdat1[8]~479 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \rfif.rdat2[7]~524 (
// Equation(s):
// rfifrdat2_7 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[7]~513_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[7]~523_combout ))))

	.dataa(\rfif.rdat2[7]~523_combout ),
	.datab(Instr_IF_20),
	.datac(\WideOr1~combout ),
	.datad(\rfif.rdat2[7]~513_combout ),
	.cin(gnd),
	.combout(rfifrdat2_7),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~524 .lut_mask = 16'hE020;
defparam \rfif.rdat2[7]~524 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \rfif.rdat1[7]~489 (
// Equation(s):
// rfifrdat1_7 = (\rfif.rdat1[7]~486_combout  & (((\rfif.rdat1[7]~488_combout ) # (!Instr_IF_21)))) # (!\rfif.rdat1[7]~486_combout  & (\rfif.rdat1[7]~481_combout  & ((Instr_IF_21))))

	.dataa(\rfif.rdat1[7]~481_combout ),
	.datab(\rfif.rdat1[7]~488_combout ),
	.datac(\rfif.rdat1[7]~486_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(rfifrdat1_7),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~489 .lut_mask = 16'hCAF0;
defparam \rfif.rdat1[7]~489 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \rfif.rdat1[7]~499 (
// Equation(s):
// rfifrdat1_71 = (Instr_IF_23 & ((\rfif.rdat1[7]~496_combout  & ((\rfif.rdat1[7]~498_combout ))) # (!\rfif.rdat1[7]~496_combout  & (\rfif.rdat1[7]~491_combout )))) # (!Instr_IF_23 & (\rfif.rdat1[7]~496_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[7]~496_combout ),
	.datac(\rfif.rdat1[7]~491_combout ),
	.datad(\rfif.rdat1[7]~498_combout ),
	.cin(gnd),
	.combout(rfifrdat1_71),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~499 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[7]~499 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \rfif.rdat2[6]~545 (
// Equation(s):
// rfifrdat2_6 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[6]~534_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[6]~544_combout )))))

	.dataa(Instr_IF_20),
	.datab(\rfif.rdat2[6]~534_combout ),
	.datac(\WideOr1~combout ),
	.datad(\rfif.rdat2[6]~544_combout ),
	.cin(gnd),
	.combout(rfifrdat2_6),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~545 .lut_mask = 16'hD080;
defparam \rfif.rdat2[6]~545 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N18
cycloneive_lcell_comb \rfif.rdat1[6]~509 (
// Equation(s):
// rfifrdat1_6 = (Instr_IF_22 & ((\rfif.rdat1[6]~506_combout  & ((\rfif.rdat1[6]~508_combout ))) # (!\rfif.rdat1[6]~506_combout  & (\rfif.rdat1[6]~501_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[6]~506_combout ))))

	.dataa(\rfif.rdat1[6]~501_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[6]~508_combout ),
	.datad(\rfif.rdat1[6]~506_combout ),
	.cin(gnd),
	.combout(rfifrdat1_6),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~509 .lut_mask = 16'hF388;
defparam \rfif.rdat1[6]~509 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N14
cycloneive_lcell_comb \rfif.rdat1[6]~519 (
// Equation(s):
// rfifrdat1_61 = (\rfif.rdat1[6]~516_combout  & (((\rfif.rdat1[6]~518_combout ) # (!Instr_IF_24)))) # (!\rfif.rdat1[6]~516_combout  & (\rfif.rdat1[6]~511_combout  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[6]~511_combout ),
	.datab(\rfif.rdat1[6]~516_combout ),
	.datac(\rfif.rdat1[6]~518_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(rfifrdat1_61),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~519 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[6]~519 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[5]~566 (
// Equation(s):
// rfifrdat2_5 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[5]~555_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[5]~565_combout )))))

	.dataa(\rfif.rdat2[5]~555_combout ),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[5]~565_combout ),
	.datad(Instr_IF_20),
	.cin(gnd),
	.combout(rfifrdat2_5),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~566 .lut_mask = 16'h88C0;
defparam \rfif.rdat2[5]~566 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[5]~529 (
// Equation(s):
// rfifrdat1_5 = (\rfif.rdat1[5]~526_combout  & ((\rfif.rdat1[5]~528_combout ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[5]~526_combout  & (((\rfif.rdat1[5]~521_combout  & Instr_IF_21))))

	.dataa(\rfif.rdat1[5]~528_combout ),
	.datab(\rfif.rdat1[5]~521_combout ),
	.datac(\rfif.rdat1[5]~526_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(rfifrdat1_5),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~529 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[5]~529 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N30
cycloneive_lcell_comb \rfif.rdat1[5]~539 (
// Equation(s):
// rfifrdat1_51 = (\rfif.rdat1[5]~536_combout  & (((\rfif.rdat1[5]~538_combout ) # (!Instr_IF_23)))) # (!\rfif.rdat1[5]~536_combout  & (\rfif.rdat1[5]~531_combout  & ((Instr_IF_23))))

	.dataa(\rfif.rdat1[5]~531_combout ),
	.datab(\rfif.rdat1[5]~538_combout ),
	.datac(\rfif.rdat1[5]~536_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(rfifrdat1_51),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~539 .lut_mask = 16'hCAF0;
defparam \rfif.rdat1[5]~539 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[4]~587 (
// Equation(s):
// rfifrdat2_4 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[4]~576_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[4]~586_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[4]~586_combout ),
	.datad(\rfif.rdat2[4]~576_combout ),
	.cin(gnd),
	.combout(rfifrdat2_4),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~587 .lut_mask = 16'hC840;
defparam \rfif.rdat2[4]~587 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \rfif.rdat1[4]~549 (
// Equation(s):
// rfifrdat1_4 = (Instr_IF_22 & ((\rfif.rdat1[4]~546_combout  & (\rfif.rdat1[4]~548_combout )) # (!\rfif.rdat1[4]~546_combout  & ((\rfif.rdat1[4]~541_combout ))))) # (!Instr_IF_22 & (\rfif.rdat1[4]~546_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[4]~546_combout ),
	.datac(\rfif.rdat1[4]~548_combout ),
	.datad(\rfif.rdat1[4]~541_combout ),
	.cin(gnd),
	.combout(rfifrdat1_4),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~549 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[4]~549 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N6
cycloneive_lcell_comb \rfif.rdat1[4]~559 (
// Equation(s):
// rfifrdat1_41 = (\rfif.rdat1[4]~556_combout  & (((\rfif.rdat1[4]~558_combout )) # (!Instr_IF_24))) # (!\rfif.rdat1[4]~556_combout  & (Instr_IF_24 & ((\rfif.rdat1[4]~551_combout ))))

	.dataa(\rfif.rdat1[4]~556_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[4]~558_combout ),
	.datad(\rfif.rdat1[4]~551_combout ),
	.cin(gnd),
	.combout(rfifrdat1_41),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~559 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[4]~559 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[3]~608 (
// Equation(s):
// rfifrdat2_3 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[3]~597_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[3]~607_combout )))))

	.dataa(\WideOr1~combout ),
	.datab(\rfif.rdat2[3]~597_combout ),
	.datac(Instr_IF_20),
	.datad(\rfif.rdat2[3]~607_combout ),
	.cin(gnd),
	.combout(rfifrdat2_3),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~608 .lut_mask = 16'h8A80;
defparam \rfif.rdat2[3]~608 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[3]~569 (
// Equation(s):
// rfifrdat1_3 = (Instr_IF_21 & ((\rfif.rdat1[3]~566_combout  & (\rfif.rdat1[3]~568_combout )) # (!\rfif.rdat1[3]~566_combout  & ((\rfif.rdat1[3]~561_combout ))))) # (!Instr_IF_21 & (((\rfif.rdat1[3]~566_combout ))))

	.dataa(\rfif.rdat1[3]~568_combout ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[3]~561_combout ),
	.datad(\rfif.rdat1[3]~566_combout ),
	.cin(gnd),
	.combout(rfifrdat1_3),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~569 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[3]~569 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[3]~579 (
// Equation(s):
// rfifrdat1_32 = (Instr_IF_23 & ((\rfif.rdat1[3]~576_combout  & ((\rfif.rdat1[3]~578_combout ))) # (!\rfif.rdat1[3]~576_combout  & (\rfif.rdat1[3]~571_combout )))) # (!Instr_IF_23 & (((\rfif.rdat1[3]~576_combout ))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[3]~571_combout ),
	.datac(\rfif.rdat1[3]~576_combout ),
	.datad(\rfif.rdat1[3]~578_combout ),
	.cin(gnd),
	.combout(rfifrdat1_32),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~579 .lut_mask = 16'hF858;
defparam \rfif.rdat1[3]~579 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N12
cycloneive_lcell_comb \rfif.rdat2[2]~629 (
// Equation(s):
// rfifrdat2_2 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[2]~618_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[2]~628_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[2]~628_combout ),
	.datad(\rfif.rdat2[2]~618_combout ),
	.cin(gnd),
	.combout(rfifrdat2_2),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~629 .lut_mask = 16'hC840;
defparam \rfif.rdat2[2]~629 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \rfif.rdat1[2]~589 (
// Equation(s):
// rfifrdat1_2 = (Instr_IF_22 & ((\rfif.rdat1[2]~586_combout  & (\rfif.rdat1[2]~588_combout )) # (!\rfif.rdat1[2]~586_combout  & ((\rfif.rdat1[2]~581_combout ))))) # (!Instr_IF_22 & (\rfif.rdat1[2]~586_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[2]~586_combout ),
	.datac(\rfif.rdat1[2]~588_combout ),
	.datad(\rfif.rdat1[2]~581_combout ),
	.cin(gnd),
	.combout(rfifrdat1_2),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~589 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[2]~589 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \rfif.rdat1[2]~599 (
// Equation(s):
// rfifrdat1_210 = (Instr_IF_24 & ((\rfif.rdat1[2]~596_combout  & (\rfif.rdat1[2]~598_combout )) # (!\rfif.rdat1[2]~596_combout  & ((\rfif.rdat1[2]~591_combout ))))) # (!Instr_IF_24 & (((\rfif.rdat1[2]~596_combout ))))

	.dataa(\rfif.rdat1[2]~598_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[2]~591_combout ),
	.datad(\rfif.rdat1[2]~596_combout ),
	.cin(gnd),
	.combout(rfifrdat1_210),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~599 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[2]~599 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[1]~650 (
// Equation(s):
// rfifrdat2_1 = (\WideOr1~combout  & ((Instr_IF_20 & (\rfif.rdat2[1]~639_combout )) # (!Instr_IF_20 & ((\rfif.rdat2[1]~649_combout )))))

	.dataa(Instr_IF_20),
	.datab(\rfif.rdat2[1]~639_combout ),
	.datac(\rfif.rdat2[1]~649_combout ),
	.datad(\WideOr1~combout ),
	.cin(gnd),
	.combout(rfifrdat2_1),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~650 .lut_mask = 16'hD800;
defparam \rfif.rdat2[1]~650 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \rfif.rdat1[1]~609 (
// Equation(s):
// rfifrdat1_1 = (\rfif.rdat1[1]~606_combout  & ((\rfif.rdat1[1]~608_combout ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[1]~606_combout  & (((\rfif.rdat1[1]~601_combout  & Instr_IF_21))))

	.dataa(\rfif.rdat1[1]~606_combout ),
	.datab(\rfif.rdat1[1]~608_combout ),
	.datac(\rfif.rdat1[1]~601_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(rfifrdat1_1),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~609 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[1]~609 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \rfif.rdat1[1]~619 (
// Equation(s):
// rfifrdat1_110 = (Instr_IF_23 & ((\rfif.rdat1[1]~616_combout  & (\rfif.rdat1[1]~618_combout )) # (!\rfif.rdat1[1]~616_combout  & ((\rfif.rdat1[1]~611_combout ))))) # (!Instr_IF_23 & (\rfif.rdat1[1]~616_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[1]~616_combout ),
	.datac(\rfif.rdat1[1]~618_combout ),
	.datad(\rfif.rdat1[1]~611_combout ),
	.cin(gnd),
	.combout(rfifrdat1_110),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~619 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[1]~619 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[0]~671 (
// Equation(s):
// rfifrdat2_0 = (\WideOr1~combout  & ((Instr_IF_20 & ((\rfif.rdat2[0]~660_combout ))) # (!Instr_IF_20 & (\rfif.rdat2[0]~670_combout ))))

	.dataa(Instr_IF_20),
	.datab(\WideOr1~combout ),
	.datac(\rfif.rdat2[0]~670_combout ),
	.datad(\rfif.rdat2[0]~660_combout ),
	.cin(gnd),
	.combout(rfifrdat2_0),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~671 .lut_mask = 16'hC840;
defparam \rfif.rdat2[0]~671 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[0]~629 (
// Equation(s):
// rfifrdat1_0 = (Instr_IF_22 & ((\rfif.rdat1[0]~626_combout  & ((\rfif.rdat1[0]~628_combout ))) # (!\rfif.rdat1[0]~626_combout  & (\rfif.rdat1[0]~621_combout )))) # (!Instr_IF_22 & (((\rfif.rdat1[0]~626_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[0]~621_combout ),
	.datac(\rfif.rdat1[0]~628_combout ),
	.datad(\rfif.rdat1[0]~626_combout ),
	.cin(gnd),
	.combout(rfifrdat1_0),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~629 .lut_mask = 16'hF588;
defparam \rfif.rdat1[0]~629 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \rfif.rdat1[0]~639 (
// Equation(s):
// rfifrdat1_01 = (Instr_IF_24 & ((\rfif.rdat1[0]~636_combout  & ((\rfif.rdat1[0]~638_combout ))) # (!\rfif.rdat1[0]~636_combout  & (\rfif.rdat1[0]~631_combout )))) # (!Instr_IF_24 & (((\rfif.rdat1[0]~636_combout ))))

	.dataa(\rfif.rdat1[0]~631_combout ),
	.datab(\rfif.rdat1[0]~638_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[0]~636_combout ),
	.cin(gnd),
	.combout(rfifrdat1_01),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~639 .lut_mask = 16'hCFA0;
defparam \rfif.rdat1[0]~639 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// \WideOr1~0_combout  = (Instr_IF_19) # ((Instr_IF_17) # ((Instr_IF_20) # (Instr_IF_18)))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_17),
	.datac(Instr_IF_20),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb WideOr1(
// Equation(s):
// \WideOr1~combout  = (\WideOr1~0_combout ) # (Instr_IF_16)

	.dataa(gnd),
	.datab(\WideOr1~0_combout ),
	.datac(Instr_IF_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr1~combout ),
	.cout());
// synopsys translate_off
defparam WideOr1.lut_mask = 16'hFCFC;
defparam WideOr1.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N30
cycloneive_lcell_comb \regs[11][31]~feeder (
// Equation(s):
// \regs[11][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (RegDst_MEM_0 & (!RegDst_MEM_2 & (RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h2000;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (!RegDst_MEM_4 & (\Decoder0~18_combout  & RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~18_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h3000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N31
dffeas \regs[11][31] (
	.clk(!CLK),
	.d(\regs[11][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][31] .is_wysiwyg = "true";
defparam \regs[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (!RegDst_MEM_0 & (!RegDst_MEM_2 & (RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'h1000;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (!RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~2_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h5000;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N25
dffeas \regs[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][31] .is_wysiwyg = "true";
defparam \regs[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[31]~11 (
// Equation(s):
// \rfif.rdat2[31]~11_combout  = (\rfif.rdat2[31]~10_combout  & ((\regs[11][31]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[31]~10_combout  & (((\regs[10][31]~q  & Instr_IF_17))))

	.dataa(\rfif.rdat2[31]~10_combout ),
	.datab(\regs[11][31]~q ),
	.datac(\regs[10][31]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~11_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~11 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[31]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (RegDst_MEM_0 & (RegDst_MEM_2 & (!RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h0800;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N2
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (!RegDst_MEM_3 & (!RegDst_MEM_4 & \Decoder0~8_combout ))

	.dataa(RegDst_MEM_3),
	.datab(RegDst_MEM_4),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h1100;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N29
dffeas \regs[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][31] .is_wysiwyg = "true";
defparam \regs[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (RegDst_MEM_0 & (RegDst_MEM_2 & (RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h8000;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (!RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~20_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h0500;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N31
dffeas \regs[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][31] .is_wysiwyg = "true";
defparam \regs[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (!RegDst_MEM_0 & (RegDst_MEM_2 & (RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h4000;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (!RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~0_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h0500;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N5
dffeas \regs[6][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][31] .is_wysiwyg = "true";
defparam \regs[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (!RegDst_MEM_0 & (RegDst_MEM_2 & (!RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h0400;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (!RegDst_MEM_3 & (\Decoder0~12_combout  & !RegDst_MEM_4))

	.dataa(gnd),
	.datab(RegDst_MEM_3),
	.datac(\Decoder0~12_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h0030;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N31
dffeas \regs[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][31] .is_wysiwyg = "true";
defparam \regs[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[31]~12 (
// Equation(s):
// \rfif.rdat2[31]~12_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[6][31]~q )) # (!Instr_IF_17 & ((\regs[4][31]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[6][31]~q ),
	.datac(\regs[4][31]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~12_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~12 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[31]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[31]~13 (
// Equation(s):
// \rfif.rdat2[31]~13_combout  = (Instr_IF_16 & ((\rfif.rdat2[31]~12_combout  & ((\regs[7][31]~q ))) # (!\rfif.rdat2[31]~12_combout  & (\regs[5][31]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[31]~12_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][31]~q ),
	.datac(\regs[7][31]~q ),
	.datad(\rfif.rdat2[31]~12_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~13_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~13 .lut_mask = 16'hF588;
defparam \rfif.rdat2[31]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \rfif.rdat2[31]~16 (
// Equation(s):
// \rfif.rdat2[31]~16_combout  = (Instr_IF_18 & (((Instr_IF_19) # (\rfif.rdat2[31]~13_combout )))) # (!Instr_IF_18 & (\rfif.rdat2[31]~15_combout  & (!Instr_IF_19)))

	.dataa(\rfif.rdat2[31]~15_combout ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[31]~13_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~16_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~16 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[31]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N16
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (RegDst_MEM_3 & (!RegDst_MEM_4 & \Decoder0~8_combout ))

	.dataa(RegDst_MEM_3),
	.datab(RegDst_MEM_4),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h2200;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N13
dffeas \regs[13][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][31] .is_wysiwyg = "true";
defparam \regs[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \regs[15][31]~feeder (
// Equation(s):
// \regs[15][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[15][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \Decoder0~39 (
// Equation(s):
// \Decoder0~39_combout  = (!RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~20_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~39 .lut_mask = 16'h5000;
defparam \Decoder0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N25
dffeas \regs[15][31] (
	.clk(!CLK),
	.d(\regs[15][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][31] .is_wysiwyg = "true";
defparam \regs[15][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \rfif.rdat2[31]~18 (
// Equation(s):
// \rfif.rdat2[31]~18_combout  = (\rfif.rdat2[31]~17_combout  & (((\regs[15][31]~q )) # (!Instr_IF_16))) # (!\rfif.rdat2[31]~17_combout  & (Instr_IF_16 & (\regs[13][31]~q )))

	.dataa(\rfif.rdat2[31]~17_combout ),
	.datab(Instr_IF_16),
	.datac(\regs[13][31]~q ),
	.datad(\regs[15][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~18_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~18 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[31]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[31]~19 (
// Equation(s):
// \rfif.rdat2[31]~19_combout  = (\rfif.rdat2[31]~16_combout  & (((\rfif.rdat2[31]~18_combout ) # (!Instr_IF_19)))) # (!\rfif.rdat2[31]~16_combout  & (\rfif.rdat2[31]~11_combout  & (Instr_IF_19)))

	.dataa(\rfif.rdat2[31]~11_combout ),
	.datab(\rfif.rdat2[31]~16_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[31]~18_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~19_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~19 .lut_mask = 16'hEC2C;
defparam \rfif.rdat2[31]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N8
cycloneive_lcell_comb \regs[27][31]~feeder (
// Equation(s):
// \regs[27][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (RegDst_MEM_4 & (\Decoder0~18_combout  & RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~18_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'hC000;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N9
dffeas \regs[27][31] (
	.clk(!CLK),
	.d(\regs[27][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][31] .is_wysiwyg = "true";
defparam \regs[27][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~20_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'hA000;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N17
dffeas \regs[31][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][31] .is_wysiwyg = "true";
defparam \regs[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N16
cycloneive_lcell_comb \rfif.rdat2[31]~8 (
// Equation(s):
// \rfif.rdat2[31]~8_combout  = (\rfif.rdat2[31]~7_combout  & (((\regs[31][31]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[31]~7_combout  & (\regs[27][31]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[31]~7_combout ),
	.datab(\regs[27][31]~q ),
	.datac(\regs[31][31]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~8_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~8 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[31]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \Decoder0~5 (
// Equation(s):
// \Decoder0~5_combout  = (\Decoder0~0_combout  & (RegDst_MEM_3 & RegDst_MEM_4))

	.dataa(\Decoder0~0_combout ),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~5 .lut_mask = 16'hA000;
defparam \Decoder0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N7
dffeas \regs[30][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][31] .is_wysiwyg = "true";
defparam \regs[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (\Decoder0~0_combout  & (!RegDst_MEM_3 & RegDst_MEM_4))

	.dataa(\Decoder0~0_combout ),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h0A00;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N5
dffeas \regs[22][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][31] .is_wysiwyg = "true";
defparam \regs[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \Decoder0~4 (
// Equation(s):
// \Decoder0~4_combout  = (RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~2_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~4 .lut_mask = 16'h0A00;
defparam \Decoder0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N7
dffeas \regs[18][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][31] .is_wysiwyg = "true";
defparam \regs[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \Decoder0~3 (
// Equation(s):
// \Decoder0~3_combout  = (RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~2_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~3 .lut_mask = 16'hA000;
defparam \Decoder0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N25
dffeas \regs[26][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][31] .is_wysiwyg = "true";
defparam \regs[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \rfif.rdat2[31]~0 (
// Equation(s):
// \rfif.rdat2[31]~0_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][31]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][31]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][31]~q ),
	.datad(\regs[26][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~0 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[31]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \rfif.rdat2[31]~1 (
// Equation(s):
// \rfif.rdat2[31]~1_combout  = (Instr_IF_18 & ((\rfif.rdat2[31]~0_combout  & (\regs[30][31]~q )) # (!\rfif.rdat2[31]~0_combout  & ((\regs[22][31]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[31]~0_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[30][31]~q ),
	.datac(\regs[22][31]~q ),
	.datad(\rfif.rdat2[31]~0_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~1 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[31]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (!RegDst_MEM_0 & (!RegDst_MEM_2 & (!RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0100;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N4
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (!RegDst_MEM_3 & (\Decoder0~14_combout  & RegDst_MEM_4))

	.dataa(RegDst_MEM_3),
	.datab(gnd),
	.datac(\Decoder0~14_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h5000;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N31
dffeas \regs[16][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][31] .is_wysiwyg = "true";
defparam \regs[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N14
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (RegDst_MEM_3 & (\Decoder0~14_combout  & RegDst_MEM_4))

	.dataa(RegDst_MEM_3),
	.datab(gnd),
	.datac(\Decoder0~14_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'hA000;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N13
dffeas \regs[24][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][31] .is_wysiwyg = "true";
defparam \regs[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[31]~4 (
// Equation(s):
// \rfif.rdat2[31]~4_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[24][31]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[16][31]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][31]~q ),
	.datad(\regs[24][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~4_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~4 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[31]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N2
cycloneive_lcell_comb \regs[28][31]~feeder (
// Equation(s):
// \regs[28][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[28][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (RegDst_MEM_3 & (\Decoder0~12_combout  & RegDst_MEM_4))

	.dataa(RegDst_MEM_3),
	.datab(gnd),
	.datac(\Decoder0~12_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'hA000;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N3
dffeas \regs[28][31] (
	.clk(!CLK),
	.d(\regs[28][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][31] .is_wysiwyg = "true";
defparam \regs[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N28
cycloneive_lcell_comb \rfif.rdat2[31]~5 (
// Equation(s):
// \rfif.rdat2[31]~5_combout  = (\rfif.rdat2[31]~4_combout  & (((\regs[28][31]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[31]~4_combout  & (\regs[20][31]~q  & (Instr_IF_18)))

	.dataa(\regs[20][31]~q ),
	.datab(\rfif.rdat2[31]~4_combout ),
	.datac(Instr_IF_18),
	.datad(\regs[28][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~5_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~5 .lut_mask = 16'hEC2C;
defparam \rfif.rdat2[31]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \rfif.rdat2[31]~6 (
// Equation(s):
// \rfif.rdat2[31]~6_combout  = (Instr_IF_16 & ((\rfif.rdat2[31]~3_combout ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((!Instr_IF_17 & \rfif.rdat2[31]~5_combout ))))

	.dataa(\rfif.rdat2[31]~3_combout ),
	.datab(Instr_IF_16),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[31]~5_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~6_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~6 .lut_mask = 16'hCBC8;
defparam \rfif.rdat2[31]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[31]~9 (
// Equation(s):
// \rfif.rdat2[31]~9_combout  = (Instr_IF_17 & ((\rfif.rdat2[31]~6_combout  & (\rfif.rdat2[31]~8_combout )) # (!\rfif.rdat2[31]~6_combout  & ((\rfif.rdat2[31]~1_combout ))))) # (!Instr_IF_17 & (((\rfif.rdat2[31]~6_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[31]~8_combout ),
	.datac(\rfif.rdat2[31]~1_combout ),
	.datad(\rfif.rdat2[31]~6_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[31]~9_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[31]~9 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[31]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \rfif.rdat1[31]~0 (
// Equation(s):
// \rfif.rdat1[31]~0_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][31]~q )) # (!Instr_IF_24 & ((\regs[18][31]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][31]~q ),
	.datad(\regs[18][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~0 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[31]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \rfif.rdat1[31]~1 (
// Equation(s):
// \rfif.rdat1[31]~1_combout  = (Instr_IF_23 & ((\rfif.rdat1[31]~0_combout  & (\regs[30][31]~q )) # (!\rfif.rdat1[31]~0_combout  & ((\regs[22][31]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[31]~0_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[31]~0_combout ),
	.datac(\regs[30][31]~q ),
	.datad(\regs[22][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~1 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[31]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \regs[23][31]~feeder (
// Equation(s):
// \regs[23][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[23][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~20_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h0A00;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N5
dffeas \regs[23][31] (
	.clk(!CLK),
	.d(\regs[23][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][31] .is_wysiwyg = "true";
defparam \regs[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \regs[19][31]~feeder (
// Equation(s):
// \regs[19][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[19][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (RegDst_MEM_4 & (\Decoder0~18_combout  & !RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~18_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h00C0;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N17
dffeas \regs[19][31] (
	.clk(!CLK),
	.d(\regs[19][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][31] .is_wysiwyg = "true";
defparam \regs[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[31]~7 (
// Equation(s):
// \rfif.rdat1[31]~7_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][31]~q )) # (!Instr_IF_23 & ((\regs[19][31]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][31]~q ),
	.datad(\regs[19][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~7_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~7 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[31]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \rfif.rdat1[31]~8 (
// Equation(s):
// \rfif.rdat1[31]~8_combout  = (Instr_IF_24 & ((\rfif.rdat1[31]~7_combout  & (\regs[31][31]~q )) # (!\rfif.rdat1[31]~7_combout  & ((\regs[27][31]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[31]~7_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[31][31]~q ),
	.datac(\regs[27][31]~q ),
	.datad(\rfif.rdat1[31]~7_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~8_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~8 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[31]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \Decoder0~6 (
// Equation(s):
// \Decoder0~6_combout  = (RegDst_MEM_0 & (!RegDst_MEM_2 & (!RegDst_MEM_1 & RegWen_MEM1)))

	.dataa(RegDst_MEM_0),
	.datab(RegDst_MEM_2),
	.datac(RegDst_MEM_1),
	.datad(RegWen_MEM),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~6 .lut_mask = 16'h0200;
defparam \Decoder0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \Decoder0~7 (
// Equation(s):
// \Decoder0~7_combout  = (RegDst_MEM_4 & (\Decoder0~6_combout  & RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~6_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~7 .lut_mask = 16'hC000;
defparam \Decoder0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \regs[25][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][31] .is_wysiwyg = "true";
defparam \regs[25][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N24
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (!RegDst_MEM_3 & (RegDst_MEM_4 & \Decoder0~8_combout ))

	.dataa(RegDst_MEM_3),
	.datab(RegDst_MEM_4),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h4400;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N5
dffeas \regs[21][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][31] .is_wysiwyg = "true";
defparam \regs[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (RegDst_MEM_4 & (\Decoder0~6_combout  & !RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~6_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h00C0;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N11
dffeas \regs[17][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][31] .is_wysiwyg = "true";
defparam \regs[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[31]~2 (
// Equation(s):
// \rfif.rdat1[31]~2_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[21][31]~q )) # (!Instr_IF_23 & ((\regs[17][31]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[21][31]~q ),
	.datad(\regs[17][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~2_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~2 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[31]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[31]~3 (
// Equation(s):
// \rfif.rdat1[31]~3_combout  = (Instr_IF_24 & ((\rfif.rdat1[31]~2_combout  & (\regs[29][31]~q )) # (!\rfif.rdat1[31]~2_combout  & ((\regs[25][31]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[31]~2_combout ))))

	.dataa(\regs[29][31]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[25][31]~q ),
	.datad(\rfif.rdat1[31]~2_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~3 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[31]~4 (
// Equation(s):
// \rfif.rdat1[31]~4_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][31]~q ))) # (!Instr_IF_24 & (\regs[16][31]~q ))))

	.dataa(\regs[16][31]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[24][31]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~4_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~4 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[31]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N30
cycloneive_lcell_comb \rfif.rdat1[31]~5 (
// Equation(s):
// \rfif.rdat1[31]~5_combout  = (\rfif.rdat1[31]~4_combout  & (((\regs[28][31]~q ) # (!Instr_IF_23)))) # (!\rfif.rdat1[31]~4_combout  & (\regs[20][31]~q  & ((Instr_IF_23))))

	.dataa(\regs[20][31]~q ),
	.datab(\regs[28][31]~q ),
	.datac(\rfif.rdat1[31]~4_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~5_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~5 .lut_mask = 16'hCAF0;
defparam \rfif.rdat1[31]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[31]~6 (
// Equation(s):
// \rfif.rdat1[31]~6_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\rfif.rdat1[31]~3_combout )) # (!Instr_IF_21 & ((\rfif.rdat1[31]~5_combout )))))

	.dataa(\rfif.rdat1[31]~3_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[31]~5_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~6_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~6 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[31]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \regs[8][31]~feeder (
// Equation(s):
// \regs[8][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][31]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~14_combout ))

	.dataa(RegDst_MEM_4),
	.datab(RegDst_MEM_3),
	.datac(gnd),
	.datad(\Decoder0~14_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h4400;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N11
dffeas \regs[8][31] (
	.clk(!CLK),
	.d(\regs[8][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][31] .is_wysiwyg = "true";
defparam \regs[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (!RegDst_MEM_4 & (\Decoder0~6_combout  & RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~6_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h3000;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N13
dffeas \regs[9][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][31] .is_wysiwyg = "true";
defparam \regs[9][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[31]~10 (
// Equation(s):
// \rfif.rdat1[31]~10_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][31]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & (\regs[8][31]~q )))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[8][31]~q ),
	.datad(\regs[9][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~10_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~10 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[31]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[31]~11 (
// Equation(s):
// \rfif.rdat1[31]~11_combout  = (\rfif.rdat1[31]~10_combout  & ((\regs[11][31]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[31]~10_combout  & (((Instr_IF_22 & \regs[10][31]~q ))))

	.dataa(\rfif.rdat1[31]~10_combout ),
	.datab(\regs[11][31]~q ),
	.datac(Instr_IF_22),
	.datad(\regs[10][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~11_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~11 .lut_mask = 16'hDA8A;
defparam \rfif.rdat1[31]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[31]~12 (
// Equation(s):
// \rfif.rdat1[31]~12_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[6][31]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[4][31]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[6][31]~q ),
	.datad(\regs[4][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~12_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~12 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[31]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[31]~13 (
// Equation(s):
// \rfif.rdat1[31]~13_combout  = (Instr_IF_21 & ((\rfif.rdat1[31]~12_combout  & (\regs[7][31]~q )) # (!\rfif.rdat1[31]~12_combout  & ((\regs[5][31]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[31]~12_combout ))))

	.dataa(\regs[7][31]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][31]~q ),
	.datad(\rfif.rdat1[31]~12_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~13_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~13 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[31]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (!RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~2_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0500;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N5
dffeas \regs[2][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][31] .is_wysiwyg = "true";
defparam \regs[2][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \regs[3][31]~feeder (
// Equation(s):
// \regs[3][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[3][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!RegDst_MEM_4 & (\Decoder0~18_combout  & !RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~18_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h0030;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N17
dffeas \regs[3][31] (
	.clk(!CLK),
	.d(\regs[3][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][31] .is_wysiwyg = "true";
defparam \regs[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[31]~15 (
// Equation(s):
// \rfif.rdat1[31]~15_combout  = (\rfif.rdat1[31]~14_combout  & (((\regs[3][31]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[31]~14_combout  & (Instr_IF_22 & (\regs[2][31]~q )))

	.dataa(\rfif.rdat1[31]~14_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[2][31]~q ),
	.datad(\regs[3][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~15_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~15 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[31]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \rfif.rdat1[31]~16 (
// Equation(s):
// \rfif.rdat1[31]~16_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\rfif.rdat1[31]~13_combout )) # (!Instr_IF_23 & ((\rfif.rdat1[31]~15_combout )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[31]~13_combout ),
	.datad(\rfif.rdat1[31]~15_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~16_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~16 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[31]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \regs[14][31]~feeder (
// Equation(s):
// \regs[14][31]~feeder_combout  = \input_a~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a),
	.cin(gnd),
	.combout(\regs[14][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][31]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (!RegDst_MEM_4 & (RegDst_MEM_3 & \Decoder0~0_combout ))

	.dataa(RegDst_MEM_4),
	.datab(gnd),
	.datac(RegDst_MEM_3),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h5000;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N21
dffeas \regs[14][31] (
	.clk(!CLK),
	.d(\regs[14][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][31] .is_wysiwyg = "true";
defparam \regs[14][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (RegDst_MEM_3 & (\Decoder0~12_combout  & !RegDst_MEM_4))

	.dataa(gnd),
	.datab(RegDst_MEM_3),
	.datac(\Decoder0~12_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'h00C0;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N23
dffeas \regs[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][31] .is_wysiwyg = "true";
defparam \regs[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[31]~17 (
// Equation(s):
// \rfif.rdat1[31]~17_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][31]~q )) # (!Instr_IF_22 & ((\regs[12][31]~q )))))

	.dataa(Instr_IF_21),
	.datab(\regs[14][31]~q ),
	.datac(Instr_IF_22),
	.datad(\regs[12][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~17_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~17 .lut_mask = 16'hE5E0;
defparam \rfif.rdat1[31]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[31]~18 (
// Equation(s):
// \rfif.rdat1[31]~18_combout  = (\rfif.rdat1[31]~17_combout  & ((\regs[15][31]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[31]~17_combout  & (((Instr_IF_21 & \regs[13][31]~q ))))

	.dataa(\rfif.rdat1[31]~17_combout ),
	.datab(\regs[15][31]~q ),
	.datac(Instr_IF_21),
	.datad(\regs[13][31]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[31]~18_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[31]~18 .lut_mask = 16'hDA8A;
defparam \rfif.rdat1[31]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \regs[27][30]~feeder (
// Equation(s):
// \regs[27][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N13
dffeas \regs[27][30] (
	.clk(!CLK),
	.d(\regs[27][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][30] .is_wysiwyg = "true";
defparam \regs[27][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[30]~27 (
// Equation(s):
// \rfif.rdat1[30]~27_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[27][30]~q ))) # (!Instr_IF_24 & (\regs[19][30]~q ))))

	.dataa(\regs[19][30]~q ),
	.datab(Instr_IF_23),
	.datac(Instr_IF_24),
	.datad(\regs[27][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~27_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~27 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[30]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \regs[31][30]~feeder (
// Equation(s):
// \regs[31][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N21
dffeas \regs[31][30] (
	.clk(!CLK),
	.d(\regs[31][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][30] .is_wysiwyg = "true";
defparam \regs[31][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \regs[23][30]~feeder (
// Equation(s):
// \regs[23][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N3
dffeas \regs[23][30] (
	.clk(!CLK),
	.d(\regs[23][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][30] .is_wysiwyg = "true";
defparam \regs[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[30]~28 (
// Equation(s):
// \rfif.rdat1[30]~28_combout  = (\rfif.rdat1[30]~27_combout  & (((\regs[31][30]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[30]~27_combout  & (Instr_IF_23 & ((\regs[23][30]~q ))))

	.dataa(\rfif.rdat1[30]~27_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[31][30]~q ),
	.datad(\regs[23][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~28_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~28 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[30]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N7
dffeas \regs[16][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][30] .is_wysiwyg = "true";
defparam \regs[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N4
cycloneive_lcell_comb \regs[20][30]~feeder (
// Equation(s):
// \regs[20][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b),
	.cin(gnd),
	.combout(\regs[20][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][30]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (!RegDst_MEM_3 & (\Decoder0~12_combout  & RegDst_MEM_4))

	.dataa(RegDst_MEM_3),
	.datab(gnd),
	.datac(\Decoder0~12_combout ),
	.datad(RegDst_MEM_4),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h5000;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N5
dffeas \regs[20][30] (
	.clk(!CLK),
	.d(\regs[20][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][30] .is_wysiwyg = "true";
defparam \regs[20][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[30]~24 (
// Equation(s):
// \rfif.rdat1[30]~24_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[20][30]~q ))) # (!Instr_IF_23 & (\regs[16][30]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[16][30]~q ),
	.datac(Instr_IF_23),
	.datad(\regs[20][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~24_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~24 .lut_mask = 16'hF4A4;
defparam \rfif.rdat1[30]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N1
dffeas \regs[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][30] .is_wysiwyg = "true";
defparam \regs[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N18
cycloneive_lcell_comb \regs[28][30]~feeder (
// Equation(s):
// \regs[28][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b),
	.cin(gnd),
	.combout(\regs[28][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][30]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N19
dffeas \regs[28][30] (
	.clk(!CLK),
	.d(\regs[28][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][30] .is_wysiwyg = "true";
defparam \regs[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[30]~25 (
// Equation(s):
// \rfif.rdat1[30]~25_combout  = (Instr_IF_24 & ((\rfif.rdat1[30]~24_combout  & ((\regs[28][30]~q ))) # (!\rfif.rdat1[30]~24_combout  & (\regs[24][30]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[30]~24_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[30]~24_combout ),
	.datac(\regs[24][30]~q ),
	.datad(\regs[28][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~25_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~25 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[30]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N3
dffeas \regs[30][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][30] .is_wysiwyg = "true";
defparam \regs[30][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \regs[26][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][30] .is_wysiwyg = "true";
defparam \regs[26][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N29
dffeas \regs[22][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][30] .is_wysiwyg = "true";
defparam \regs[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[30]~22 (
// Equation(s):
// \rfif.rdat1[30]~22_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][30]~q ))) # (!Instr_IF_23 & (\regs[18][30]~q ))))

	.dataa(\regs[18][30]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[22][30]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~22_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~22 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[30]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[30]~23 (
// Equation(s):
// \rfif.rdat1[30]~23_combout  = (Instr_IF_24 & ((\rfif.rdat1[30]~22_combout  & (\regs[30][30]~q )) # (!\rfif.rdat1[30]~22_combout  & ((\regs[26][30]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[30]~22_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[30][30]~q ),
	.datac(\regs[26][30]~q ),
	.datad(\rfif.rdat1[30]~22_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~23_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~23 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[30]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[30]~26 (
// Equation(s):
// \rfif.rdat1[30]~26_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[30]~23_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[30]~25_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[30]~25_combout ),
	.datad(\rfif.rdat1[30]~23_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~26_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~26 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[30]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N29
dffeas \regs[21][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][30] .is_wysiwyg = "true";
defparam \regs[21][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N10
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (RegDst_MEM_3 & (RegDst_MEM_4 & \Decoder0~8_combout ))

	.dataa(RegDst_MEM_3),
	.datab(RegDst_MEM_4),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h8800;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N11
dffeas \regs[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][30] .is_wysiwyg = "true";
defparam \regs[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N19
dffeas \regs[17][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][30] .is_wysiwyg = "true";
defparam \regs[17][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \regs[25][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][30] .is_wysiwyg = "true";
defparam \regs[25][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[30]~20 (
// Equation(s):
// \rfif.rdat1[30]~20_combout  = (Instr_IF_24 & (((\regs[25][30]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][30]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][30]~q ),
	.datac(\regs[25][30]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~20_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~20 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[30]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[30]~21 (
// Equation(s):
// \rfif.rdat1[30]~21_combout  = (Instr_IF_23 & ((\rfif.rdat1[30]~20_combout  & ((\regs[29][30]~q ))) # (!\rfif.rdat1[30]~20_combout  & (\regs[21][30]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[30]~20_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[21][30]~q ),
	.datac(\regs[29][30]~q ),
	.datad(\rfif.rdat1[30]~20_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~21_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~21 .lut_mask = 16'hF588;
defparam \rfif.rdat1[30]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N25
dffeas \regs[2][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][30] .is_wysiwyg = "true";
defparam \regs[2][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[30]~34 (
// Equation(s):
// \rfif.rdat1[30]~34_combout  = (Instr_IF_22 & (((\regs[2][30]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[0][30]~q  & ((!Instr_IF_21))))

	.dataa(\regs[0][30]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[2][30]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~34_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~34 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[30]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!RegDst_MEM_4 & (\Decoder0~6_combout  & !RegDst_MEM_3))

	.dataa(gnd),
	.datab(RegDst_MEM_4),
	.datac(\Decoder0~6_combout ),
	.datad(RegDst_MEM_3),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h0030;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N19
dffeas \regs[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][30] .is_wysiwyg = "true";
defparam \regs[1][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N29
dffeas \regs[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][30] .is_wysiwyg = "true";
defparam \regs[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[30]~35 (
// Equation(s):
// \rfif.rdat1[30]~35_combout  = (Instr_IF_21 & ((\rfif.rdat1[30]~34_combout  & ((\regs[3][30]~q ))) # (!\rfif.rdat1[30]~34_combout  & (\regs[1][30]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[30]~34_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[30]~34_combout ),
	.datac(\regs[1][30]~q ),
	.datad(\regs[3][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~35_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~35 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[30]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N9
dffeas \regs[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][30] .is_wysiwyg = "true";
defparam \regs[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N27
dffeas \regs[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][30] .is_wysiwyg = "true";
defparam \regs[9][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N13
dffeas \regs[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][30] .is_wysiwyg = "true";
defparam \regs[10][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N19
dffeas \regs[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][30] .is_wysiwyg = "true";
defparam \regs[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[30]~32 (
// Equation(s):
// \rfif.rdat1[30]~32_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][30]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][30]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][30]~q ),
	.datad(\regs[8][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~32_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~32 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[30]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[30]~33 (
// Equation(s):
// \rfif.rdat1[30]~33_combout  = (Instr_IF_21 & ((\rfif.rdat1[30]~32_combout  & (\regs[11][30]~q )) # (!\rfif.rdat1[30]~32_combout  & ((\regs[9][30]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[30]~32_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][30]~q ),
	.datac(\regs[9][30]~q ),
	.datad(\rfif.rdat1[30]~32_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~33_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~33 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[30]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[30]~36 (
// Equation(s):
// \rfif.rdat1[30]~36_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[30]~33_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[30]~35_combout ))))

	.dataa(\rfif.rdat1[30]~35_combout ),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[30]~33_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~36_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~36 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[30]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N31
dffeas \regs[15][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][30] .is_wysiwyg = "true";
defparam \regs[15][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \regs[13][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][30] .is_wysiwyg = "true";
defparam \regs[13][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \rfif.rdat1[30]~37 (
// Equation(s):
// \rfif.rdat1[30]~37_combout  = (Instr_IF_21 & (((\regs[13][30]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][30]~q  & ((!Instr_IF_22))))

	.dataa(\regs[12][30]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][30]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~37_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~37 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[30]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N9
dffeas \regs[14][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][30] .is_wysiwyg = "true";
defparam \regs[14][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \rfif.rdat1[30]~38 (
// Equation(s):
// \rfif.rdat1[30]~38_combout  = (Instr_IF_22 & ((\rfif.rdat1[30]~37_combout  & (\regs[15][30]~q )) # (!\rfif.rdat1[30]~37_combout  & ((\regs[14][30]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[30]~37_combout ))))

	.dataa(\regs[15][30]~q ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[30]~37_combout ),
	.datad(\regs[14][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~38_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~38 .lut_mask = 16'hBCB0;
defparam \rfif.rdat1[30]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \regs[5][30]~feeder (
// Equation(s):
// \regs[5][30]~feeder_combout  = \input_b~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[5][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][30]~feeder .lut_mask = 16'hF0F0;
defparam \regs[5][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N5
dffeas \regs[5][30] (
	.clk(!CLK),
	.d(\regs[5][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][30] .is_wysiwyg = "true";
defparam \regs[5][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N31
dffeas \regs[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][30] .is_wysiwyg = "true";
defparam \regs[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \rfif.rdat1[30]~30 (
// Equation(s):
// \rfif.rdat1[30]~30_combout  = (Instr_IF_21 & ((\regs[5][30]~q ) # ((Instr_IF_22)))) # (!Instr_IF_21 & (((!Instr_IF_22 & \regs[4][30]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[5][30]~q ),
	.datac(Instr_IF_22),
	.datad(\regs[4][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~30 .lut_mask = 16'hADA8;
defparam \rfif.rdat1[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N25
dffeas \regs[7][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][30] .is_wysiwyg = "true";
defparam \regs[7][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N9
dffeas \regs[6][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][30] .is_wysiwyg = "true";
defparam \regs[6][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[30]~31 (
// Equation(s):
// \rfif.rdat1[30]~31_combout  = (\rfif.rdat1[30]~30_combout  & (((\regs[7][30]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[30]~30_combout  & (Instr_IF_22 & ((\regs[6][30]~q ))))

	.dataa(\rfif.rdat1[30]~30_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[7][30]~q ),
	.datad(\regs[6][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[30]~31_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[30]~31 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[30]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[30]~33 (
// Equation(s):
// \rfif.rdat2[30]~33_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][30]~q ))) # (!Instr_IF_17 & (\regs[8][30]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][30]~q ),
	.datad(\regs[10][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~33_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~33 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N8
cycloneive_lcell_comb \rfif.rdat2[30]~34 (
// Equation(s):
// \rfif.rdat2[30]~34_combout  = (Instr_IF_16 & ((\rfif.rdat2[30]~33_combout  & ((\regs[11][30]~q ))) # (!\rfif.rdat2[30]~33_combout  & (\regs[9][30]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[30]~33_combout ))))

	.dataa(\regs[9][30]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[11][30]~q ),
	.datad(\rfif.rdat2[30]~33_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~34_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~34 .lut_mask = 16'hF388;
defparam \rfif.rdat2[30]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!RegDst_MEM_4 & (!RegDst_MEM_3 & \Decoder0~14_combout ))

	.dataa(RegDst_MEM_4),
	.datab(RegDst_MEM_3),
	.datac(\Decoder0~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h1010;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N31
dffeas \regs[0][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][30] .is_wysiwyg = "true";
defparam \regs[0][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[30]~35 (
// Equation(s):
// \rfif.rdat2[30]~35_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[2][30]~q ))) # (!Instr_IF_17 & (\regs[0][30]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][30]~q ),
	.datad(\regs[2][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~35_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~35 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[30]~36 (
// Equation(s):
// \rfif.rdat2[30]~36_combout  = (Instr_IF_16 & ((\rfif.rdat2[30]~35_combout  & (\regs[3][30]~q )) # (!\rfif.rdat2[30]~35_combout  & ((\regs[1][30]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[30]~35_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[30]~35_combout ),
	.datac(\regs[3][30]~q ),
	.datad(\regs[1][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~36_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~36 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[30]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \rfif.rdat2[30]~37 (
// Equation(s):
// \rfif.rdat2[30]~37_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[30]~34_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[30]~36_combout )))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[30]~34_combout ),
	.datac(\rfif.rdat2[30]~36_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~37_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~37 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[30]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \rfif.rdat2[30]~39 (
// Equation(s):
// \rfif.rdat2[30]~39_combout  = (\rfif.rdat2[30]~38_combout  & ((\regs[15][30]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[30]~38_combout  & (((\regs[14][30]~q  & Instr_IF_17))))

	.dataa(\rfif.rdat2[30]~38_combout ),
	.datab(\regs[15][30]~q ),
	.datac(\regs[14][30]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~39_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~39 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[30]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[30]~31 (
// Equation(s):
// \rfif.rdat2[30]~31_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][30]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][30]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][30]~q ),
	.datad(\regs[5][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~31_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~31 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[30]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[30]~32 (
// Equation(s):
// \rfif.rdat2[30]~32_combout  = (Instr_IF_17 & ((\rfif.rdat2[30]~31_combout  & (\regs[7][30]~q )) # (!\rfif.rdat2[30]~31_combout  & ((\regs[6][30]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[30]~31_combout ))))

	.dataa(\regs[7][30]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[6][30]~q ),
	.datad(\rfif.rdat2[30]~31_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~32_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~32 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[30]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \rfif.rdat2[30]~40 (
// Equation(s):
// \rfif.rdat2[30]~40_combout  = (Instr_IF_18 & ((\rfif.rdat2[30]~37_combout  & (\rfif.rdat2[30]~39_combout )) # (!\rfif.rdat2[30]~37_combout  & ((\rfif.rdat2[30]~32_combout ))))) # (!Instr_IF_18 & (\rfif.rdat2[30]~37_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[30]~37_combout ),
	.datac(\rfif.rdat2[30]~39_combout ),
	.datad(\rfif.rdat2[30]~32_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~40_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~40 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[30]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[30]~21 (
// Equation(s):
// \rfif.rdat2[30]~21_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][30]~q ))) # (!Instr_IF_19 & (\regs[17][30]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][30]~q ),
	.datad(\regs[25][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~21_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~21 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \rfif.rdat2[30]~22 (
// Equation(s):
// \rfif.rdat2[30]~22_combout  = (Instr_IF_18 & ((\rfif.rdat2[30]~21_combout  & ((\regs[29][30]~q ))) # (!\rfif.rdat2[30]~21_combout  & (\regs[21][30]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[30]~21_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[30]~21_combout ),
	.datac(\regs[21][30]~q ),
	.datad(\regs[29][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~22_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~22 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[30]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[30]~25 (
// Equation(s):
// \rfif.rdat2[30]~25_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][30]~q ))) # (!Instr_IF_18 & (\regs[16][30]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][30]~q ),
	.datad(\regs[20][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~25_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~25 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[30]~26 (
// Equation(s):
// \rfif.rdat2[30]~26_combout  = (Instr_IF_19 & ((\rfif.rdat2[30]~25_combout  & ((\regs[28][30]~q ))) # (!\rfif.rdat2[30]~25_combout  & (\regs[24][30]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[30]~25_combout ))))

	.dataa(\regs[24][30]~q ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[30]~25_combout ),
	.datad(\regs[28][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~26_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~26 .lut_mask = 16'hF838;
defparam \rfif.rdat2[30]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N31
dffeas \regs[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][30] .is_wysiwyg = "true";
defparam \regs[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \rfif.rdat2[30]~23 (
// Equation(s):
// \rfif.rdat2[30]~23_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][30]~q ))) # (!Instr_IF_18 & (\regs[18][30]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][30]~q ),
	.datad(\regs[22][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~23_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~23 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[30]~24 (
// Equation(s):
// \rfif.rdat2[30]~24_combout  = (Instr_IF_19 & ((\rfif.rdat2[30]~23_combout  & ((\regs[30][30]~q ))) # (!\rfif.rdat2[30]~23_combout  & (\regs[26][30]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[30]~23_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][30]~q ),
	.datac(\regs[30][30]~q ),
	.datad(\rfif.rdat2[30]~23_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~24_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~24 .lut_mask = 16'hF588;
defparam \rfif.rdat2[30]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[30]~27 (
// Equation(s):
// \rfif.rdat2[30]~27_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[30]~24_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[30]~26_combout ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[30]~26_combout ),
	.datad(\rfif.rdat2[30]~24_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~27_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~27 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[30]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[30]~29 (
// Equation(s):
// \rfif.rdat2[30]~29_combout  = (\rfif.rdat2[30]~28_combout  & (((\regs[31][30]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[30]~28_combout  & (Instr_IF_18 & (\regs[23][30]~q )))

	.dataa(\rfif.rdat2[30]~28_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[23][30]~q ),
	.datad(\regs[31][30]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~29_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~29 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[30]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[30]~30 (
// Equation(s):
// \rfif.rdat2[30]~30_combout  = (Instr_IF_16 & ((\rfif.rdat2[30]~27_combout  & ((\rfif.rdat2[30]~29_combout ))) # (!\rfif.rdat2[30]~27_combout  & (\rfif.rdat2[30]~22_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[30]~27_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[30]~22_combout ),
	.datac(\rfif.rdat2[30]~27_combout ),
	.datad(\rfif.rdat2[30]~29_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[30]~30 .lut_mask = 16'hF858;
defparam \rfif.rdat2[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N25
dffeas \regs[26][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][29] .is_wysiwyg = "true";
defparam \regs[26][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N3
dffeas \regs[18][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][29] .is_wysiwyg = "true";
defparam \regs[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[29]~40 (
// Equation(s):
// \rfif.rdat1[29]~40_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][29]~q )) # (!Instr_IF_24 & ((\regs[18][29]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][29]~q ),
	.datad(\regs[18][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~40_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~40 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[29]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N29
dffeas \regs[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][29] .is_wysiwyg = "true";
defparam \regs[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \regs[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][29] .is_wysiwyg = "true";
defparam \regs[22][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[29]~41 (
// Equation(s):
// \rfif.rdat1[29]~41_combout  = (Instr_IF_23 & ((\rfif.rdat1[29]~40_combout  & (\regs[30][29]~q )) # (!\rfif.rdat1[29]~40_combout  & ((\regs[22][29]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[29]~40_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[29]~40_combout ),
	.datac(\regs[30][29]~q ),
	.datad(\regs[22][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~41_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~41 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[29]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N29
dffeas \regs[25][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][29] .is_wysiwyg = "true";
defparam \regs[25][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \regs[29][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][29] .is_wysiwyg = "true";
defparam \regs[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[29]~43 (
// Equation(s):
// \rfif.rdat1[29]~43_combout  = (\rfif.rdat1[29]~42_combout  & (((\regs[29][29]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[29]~42_combout  & (Instr_IF_24 & (\regs[25][29]~q )))

	.dataa(\rfif.rdat1[29]~42_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[25][29]~q ),
	.datad(\regs[29][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~43_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~43 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[29]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N11
dffeas \regs[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][29] .is_wysiwyg = "true";
defparam \regs[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N25
dffeas \regs[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][29] .is_wysiwyg = "true";
defparam \regs[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N10
cycloneive_lcell_comb \rfif.rdat1[29]~44 (
// Equation(s):
// \rfif.rdat1[29]~44_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[24][29]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[16][29]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[24][29]~q ),
	.datad(\regs[16][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~44_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~44 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[29]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N0
cycloneive_lcell_comb \regs[20][29]~feeder (
// Equation(s):
// \regs[20][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N1
dffeas \regs[20][29] (
	.clk(!CLK),
	.d(\regs[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][29] .is_wysiwyg = "true";
defparam \regs[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[29]~45 (
// Equation(s):
// \rfif.rdat1[29]~45_combout  = (Instr_IF_23 & ((\rfif.rdat1[29]~44_combout  & (\regs[28][29]~q )) # (!\rfif.rdat1[29]~44_combout  & ((\regs[20][29]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[29]~44_combout ))))

	.dataa(\regs[28][29]~q ),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[29]~44_combout ),
	.datad(\regs[20][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~45_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~45 .lut_mask = 16'hBCB0;
defparam \rfif.rdat1[29]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \rfif.rdat1[29]~46 (
// Equation(s):
// \rfif.rdat1[29]~46_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\rfif.rdat1[29]~43_combout )) # (!Instr_IF_21 & ((\rfif.rdat1[29]~45_combout )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[29]~43_combout ),
	.datad(\rfif.rdat1[29]~45_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~46_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~46 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[29]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \regs[31][29]~feeder (
// Equation(s):
// \regs[31][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[31][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N25
dffeas \regs[31][29] (
	.clk(!CLK),
	.d(\regs[31][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][29] .is_wysiwyg = "true";
defparam \regs[31][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \regs[23][29]~feeder (
// Equation(s):
// \regs[23][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N27
dffeas \regs[23][29] (
	.clk(!CLK),
	.d(\regs[23][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][29] .is_wysiwyg = "true";
defparam \regs[23][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \regs[19][29]~feeder (
// Equation(s):
// \regs[19][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[19][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N9
dffeas \regs[19][29] (
	.clk(!CLK),
	.d(\regs[19][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][29] .is_wysiwyg = "true";
defparam \regs[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \rfif.rdat1[29]~47 (
// Equation(s):
// \rfif.rdat1[29]~47_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][29]~q )) # (!Instr_IF_23 & ((\regs[19][29]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][29]~q ),
	.datad(\regs[19][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~47_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~47 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[29]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \regs[27][29]~feeder (
// Equation(s):
// \regs[27][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[27][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N29
dffeas \regs[27][29] (
	.clk(!CLK),
	.d(\regs[27][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][29] .is_wysiwyg = "true";
defparam \regs[27][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \rfif.rdat1[29]~48 (
// Equation(s):
// \rfif.rdat1[29]~48_combout  = (Instr_IF_24 & ((\rfif.rdat1[29]~47_combout  & (\regs[31][29]~q )) # (!\rfif.rdat1[29]~47_combout  & ((\regs[27][29]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[29]~47_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[31][29]~q ),
	.datac(\rfif.rdat1[29]~47_combout ),
	.datad(\regs[27][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~48_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~48 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[29]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N0
cycloneive_lcell_comb \regs[14][29]~feeder (
// Equation(s):
// \regs[14][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N1
dffeas \regs[14][29] (
	.clk(!CLK),
	.d(\regs[14][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][29] .is_wysiwyg = "true";
defparam \regs[14][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \rfif.rdat1[29]~57 (
// Equation(s):
// \rfif.rdat1[29]~57_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[14][29]~q ))) # (!Instr_IF_22 & (\regs[12][29]~q ))))

	.dataa(\regs[12][29]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[14][29]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~57_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~57 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[29]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N21
dffeas \regs[15][29] (
	.clk(!CLK),
	.d(input_b1),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][29] .is_wysiwyg = "true";
defparam \regs[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N17
dffeas \regs[13][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][29] .is_wysiwyg = "true";
defparam \regs[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[29]~58 (
// Equation(s):
// \rfif.rdat1[29]~58_combout  = (\rfif.rdat1[29]~57_combout  & ((\regs[15][29]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[29]~57_combout  & (((\regs[13][29]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[29]~57_combout ),
	.datab(\regs[15][29]~q ),
	.datac(\regs[13][29]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~58_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~58 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[29]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \regs[6][29]~feeder (
// Equation(s):
// \regs[6][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N9
dffeas \regs[6][29] (
	.clk(!CLK),
	.d(\regs[6][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][29] .is_wysiwyg = "true";
defparam \regs[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \rfif.rdat1[29]~52 (
// Equation(s):
// \rfif.rdat1[29]~52_combout  = (Instr_IF_22 & (((\regs[6][29]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[4][29]~q  & ((!Instr_IF_21))))

	.dataa(\regs[4][29]~q ),
	.datab(\regs[6][29]~q ),
	.datac(Instr_IF_22),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~52_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~52 .lut_mask = 16'hF0CA;
defparam \rfif.rdat1[29]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \regs[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][29] .is_wysiwyg = "true";
defparam \regs[5][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N19
dffeas \regs[7][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][29] .is_wysiwyg = "true";
defparam \regs[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[29]~53 (
// Equation(s):
// \rfif.rdat1[29]~53_combout  = (Instr_IF_21 & ((\rfif.rdat1[29]~52_combout  & ((\regs[7][29]~q ))) # (!\rfif.rdat1[29]~52_combout  & (\regs[5][29]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[29]~52_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[29]~52_combout ),
	.datac(\regs[5][29]~q ),
	.datad(\regs[7][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~53_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~53 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[29]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N17
dffeas \regs[2][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][29] .is_wysiwyg = "true";
defparam \regs[2][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \regs[1][29]~feeder (
// Equation(s):
// \regs[1][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[1][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][29]~feeder .lut_mask = 16'hF0F0;
defparam \regs[1][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N21
dffeas \regs[1][29] (
	.clk(!CLK),
	.d(\regs[1][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][29] .is_wysiwyg = "true";
defparam \regs[1][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N19
dffeas \regs[0][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][29] .is_wysiwyg = "true";
defparam \regs[0][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \rfif.rdat1[29]~54 (
// Equation(s):
// \rfif.rdat1[29]~54_combout  = (Instr_IF_21 & ((\regs[1][29]~q ) # ((Instr_IF_22)))) # (!Instr_IF_21 & (((\regs[0][29]~q  & !Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[1][29]~q ),
	.datac(\regs[0][29]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~54_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~54 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[29]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[29]~55 (
// Equation(s):
// \rfif.rdat1[29]~55_combout  = (Instr_IF_22 & ((\rfif.rdat1[29]~54_combout  & (\regs[3][29]~q )) # (!\rfif.rdat1[29]~54_combout  & ((\regs[2][29]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[29]~54_combout ))))

	.dataa(\regs[3][29]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[2][29]~q ),
	.datad(\rfif.rdat1[29]~54_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~55_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~55 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[29]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[29]~56 (
// Equation(s):
// \rfif.rdat1[29]~56_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & (\rfif.rdat1[29]~53_combout )) # (!Instr_IF_23 & ((\rfif.rdat1[29]~55_combout )))))

	.dataa(\rfif.rdat1[29]~53_combout ),
	.datab(\rfif.rdat1[29]~55_combout ),
	.datac(Instr_IF_24),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~56_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~56 .lut_mask = 16'hFA0C;
defparam \rfif.rdat1[29]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \regs[8][29]~feeder (
// Equation(s):
// \regs[8][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[8][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[8][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N13
dffeas \regs[8][29] (
	.clk(!CLK),
	.d(\regs[8][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][29] .is_wysiwyg = "true";
defparam \regs[8][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N11
dffeas \regs[9][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][29] .is_wysiwyg = "true";
defparam \regs[9][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[29]~50 (
// Equation(s):
// \rfif.rdat1[29]~50_combout  = (Instr_IF_21 & (((\regs[9][29]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[8][29]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[8][29]~q ),
	.datac(\regs[9][29]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~50_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~50 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[29]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N1
dffeas \regs[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][29] .is_wysiwyg = "true";
defparam \regs[11][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \regs[10][29]~feeder (
// Equation(s):
// \regs[10][29]~feeder_combout  = \input_b~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b1),
	.cin(gnd),
	.combout(\regs[10][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][29]~feeder .lut_mask = 16'hFF00;
defparam \regs[10][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N7
dffeas \regs[10][29] (
	.clk(!CLK),
	.d(\regs[10][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][29] .is_wysiwyg = "true";
defparam \regs[10][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[29]~51 (
// Equation(s):
// \rfif.rdat1[29]~51_combout  = (\rfif.rdat1[29]~50_combout  & (((\regs[11][29]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[29]~50_combout  & (Instr_IF_22 & ((\regs[10][29]~q ))))

	.dataa(\rfif.rdat1[29]~50_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[11][29]~q ),
	.datad(\regs[10][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[29]~51_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[29]~51 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[29]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[29]~52 (
// Equation(s):
// \rfif.rdat2[29]~52_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[9][29]~q )) # (!Instr_IF_16 & ((\regs[8][29]~q )))))

	.dataa(\regs[9][29]~q ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\regs[8][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~52_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~52 .lut_mask = 16'hE3E0;
defparam \rfif.rdat2[29]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[29]~53 (
// Equation(s):
// \rfif.rdat2[29]~53_combout  = (Instr_IF_17 & ((\rfif.rdat2[29]~52_combout  & (\regs[11][29]~q )) # (!\rfif.rdat2[29]~52_combout  & ((\regs[10][29]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[29]~52_combout ))))

	.dataa(\regs[11][29]~q ),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[29]~52_combout ),
	.datad(\regs[10][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~53_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~53 .lut_mask = 16'hBCB0;
defparam \rfif.rdat2[29]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N7
dffeas \regs[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][29] .is_wysiwyg = "true";
defparam \regs[4][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[29]~54 (
// Equation(s):
// \rfif.rdat2[29]~54_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[6][29]~q )) # (!Instr_IF_17 & ((\regs[4][29]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[6][29]~q ),
	.datac(\regs[4][29]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~54_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~54 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[29]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[29]~55 (
// Equation(s):
// \rfif.rdat2[29]~55_combout  = (Instr_IF_16 & ((\rfif.rdat2[29]~54_combout  & (\regs[7][29]~q )) # (!\rfif.rdat2[29]~54_combout  & ((\regs[5][29]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[29]~54_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[29]~54_combout ),
	.datac(\regs[7][29]~q ),
	.datad(\regs[5][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~55_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~55 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[29]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \rfif.rdat2[29]~58 (
// Equation(s):
// \rfif.rdat2[29]~58_combout  = (Instr_IF_18 & (((\rfif.rdat2[29]~55_combout ) # (Instr_IF_19)))) # (!Instr_IF_18 & (\rfif.rdat2[29]~57_combout  & ((!Instr_IF_19))))

	.dataa(\rfif.rdat2[29]~57_combout ),
	.datab(\rfif.rdat2[29]~55_combout ),
	.datac(Instr_IF_18),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~58_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~58 .lut_mask = 16'hF0CA;
defparam \rfif.rdat2[29]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \rfif.rdat2[29]~60 (
// Equation(s):
// \rfif.rdat2[29]~60_combout  = (\rfif.rdat2[29]~59_combout  & (((\regs[15][29]~q )) # (!Instr_IF_16))) # (!\rfif.rdat2[29]~59_combout  & (Instr_IF_16 & (\regs[13][29]~q )))

	.dataa(\rfif.rdat2[29]~59_combout ),
	.datab(Instr_IF_16),
	.datac(\regs[13][29]~q ),
	.datad(\regs[15][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~60_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~60 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[29]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \rfif.rdat2[29]~61 (
// Equation(s):
// \rfif.rdat2[29]~61_combout  = (Instr_IF_19 & ((\rfif.rdat2[29]~58_combout  & ((\rfif.rdat2[29]~60_combout ))) # (!\rfif.rdat2[29]~58_combout  & (\rfif.rdat2[29]~53_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[29]~58_combout ))))

	.dataa(\rfif.rdat2[29]~53_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[29]~58_combout ),
	.datad(\rfif.rdat2[29]~60_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~61_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~61 .lut_mask = 16'hF838;
defparam \rfif.rdat2[29]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \rfif.rdat2[29]~42 (
// Equation(s):
// \rfif.rdat2[29]~42_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][29]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][29]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][29]~q ),
	.datad(\regs[26][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~42_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~42 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[29]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \rfif.rdat2[29]~43 (
// Equation(s):
// \rfif.rdat2[29]~43_combout  = (Instr_IF_18 & ((\rfif.rdat2[29]~42_combout  & (\regs[30][29]~q )) # (!\rfif.rdat2[29]~42_combout  & ((\regs[22][29]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[29]~42_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[30][29]~q ),
	.datac(\regs[22][29]~q ),
	.datad(\rfif.rdat2[29]~42_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~43_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~43 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[29]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[29]~49 (
// Equation(s):
// \rfif.rdat2[29]~49_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[23][29]~q )) # (!Instr_IF_18 & ((\regs[19][29]~q )))))

	.dataa(\regs[23][29]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[19][29]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~49_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~49 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[29]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \rfif.rdat2[29]~50 (
// Equation(s):
// \rfif.rdat2[29]~50_combout  = (\rfif.rdat2[29]~49_combout  & (((\regs[31][29]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[29]~49_combout  & (\regs[27][29]~q  & ((Instr_IF_19))))

	.dataa(\regs[27][29]~q ),
	.datab(\regs[31][29]~q ),
	.datac(\rfif.rdat2[29]~49_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~50_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~50 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[29]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[29]~45 (
// Equation(s):
// \rfif.rdat2[29]~45_combout  = (\rfif.rdat2[29]~44_combout  & (((\regs[29][29]~q )) # (!Instr_IF_19))) # (!\rfif.rdat2[29]~44_combout  & (Instr_IF_19 & ((\regs[25][29]~q ))))

	.dataa(\rfif.rdat2[29]~44_combout ),
	.datab(Instr_IF_19),
	.datac(\regs[29][29]~q ),
	.datad(\regs[25][29]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~45_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~45 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[29]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[29]~48 (
// Equation(s):
// \rfif.rdat2[29]~48_combout  = (Instr_IF_16 & (((\rfif.rdat2[29]~45_combout ) # (Instr_IF_17)))) # (!Instr_IF_16 & (\rfif.rdat2[29]~47_combout  & ((!Instr_IF_17))))

	.dataa(\rfif.rdat2[29]~47_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[29]~45_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~48_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~48 .lut_mask = 16'hCCE2;
defparam \rfif.rdat2[29]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[29]~51 (
// Equation(s):
// \rfif.rdat2[29]~51_combout  = (\rfif.rdat2[29]~48_combout  & (((\rfif.rdat2[29]~50_combout ) # (!Instr_IF_17)))) # (!\rfif.rdat2[29]~48_combout  & (\rfif.rdat2[29]~43_combout  & ((Instr_IF_17))))

	.dataa(\rfif.rdat2[29]~43_combout ),
	.datab(\rfif.rdat2[29]~50_combout ),
	.datac(\rfif.rdat2[29]~48_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[29]~51_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[29]~51 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[29]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N22
cycloneive_lcell_comb \regs[24][28]~feeder (
// Equation(s):
// \regs[24][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N23
dffeas \regs[24][28] (
	.clk(!CLK),
	.d(\regs[24][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][28] .is_wysiwyg = "true";
defparam \regs[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N7
dffeas \regs[28][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][28] .is_wysiwyg = "true";
defparam \regs[28][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N22
cycloneive_lcell_comb \regs[20][28]~feeder (
// Equation(s):
// \regs[20][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N23
dffeas \regs[20][28] (
	.clk(!CLK),
	.d(\regs[20][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][28] .is_wysiwyg = "true";
defparam \regs[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N17
dffeas \regs[16][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][28] .is_wysiwyg = "true";
defparam \regs[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[28]~64 (
// Equation(s):
// \rfif.rdat1[28]~64_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[20][28]~q )) # (!Instr_IF_23 & ((\regs[16][28]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[20][28]~q ),
	.datad(\regs[16][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~64_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~64 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[28]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[28]~65 (
// Equation(s):
// \rfif.rdat1[28]~65_combout  = (Instr_IF_24 & ((\rfif.rdat1[28]~64_combout  & ((\regs[28][28]~q ))) # (!\rfif.rdat1[28]~64_combout  & (\regs[24][28]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[28]~64_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[24][28]~q ),
	.datac(\regs[28][28]~q ),
	.datad(\rfif.rdat1[28]~64_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~65_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~65 .lut_mask = 16'hF588;
defparam \rfif.rdat1[28]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N13
dffeas \regs[22][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][28] .is_wysiwyg = "true";
defparam \regs[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \rfif.rdat1[28]~62 (
// Equation(s):
// \rfif.rdat1[28]~62_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][28]~q ))) # (!Instr_IF_23 & (\regs[18][28]~q ))))

	.dataa(\regs[18][28]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[22][28]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~62_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~62 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[28]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N1
dffeas \regs[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][28] .is_wysiwyg = "true";
defparam \regs[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N7
dffeas \regs[30][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][28] .is_wysiwyg = "true";
defparam \regs[30][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[28]~63 (
// Equation(s):
// \rfif.rdat1[28]~63_combout  = (Instr_IF_24 & ((\rfif.rdat1[28]~62_combout  & ((\regs[30][28]~q ))) # (!\rfif.rdat1[28]~62_combout  & (\regs[26][28]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[28]~62_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[28]~62_combout ),
	.datac(\regs[26][28]~q ),
	.datad(\regs[30][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~63_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~63 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[28]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[28]~66 (
// Equation(s):
// \rfif.rdat1[28]~66_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[28]~63_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[28]~65_combout ))))

	.dataa(\rfif.rdat1[28]~65_combout ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[28]~63_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~66_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~66 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[28]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \regs[31][28]~feeder (
// Equation(s):
// \regs[31][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N1
dffeas \regs[31][28] (
	.clk(!CLK),
	.d(\regs[31][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][28] .is_wysiwyg = "true";
defparam \regs[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \regs[23][28]~feeder (
// Equation(s):
// \regs[23][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N23
dffeas \regs[23][28] (
	.clk(!CLK),
	.d(\regs[23][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][28] .is_wysiwyg = "true";
defparam \regs[23][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \regs[27][28]~feeder (
// Equation(s):
// \regs[27][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b2),
	.cin(gnd),
	.combout(\regs[27][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][28]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N9
dffeas \regs[27][28] (
	.clk(!CLK),
	.d(\regs[27][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][28] .is_wysiwyg = "true";
defparam \regs[27][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \regs[19][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][28] .is_wysiwyg = "true";
defparam \regs[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \rfif.rdat1[28]~67 (
// Equation(s):
// \rfif.rdat1[28]~67_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][28]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][28]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][28]~q ),
	.datad(\regs[19][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~67_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~67 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[28]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[28]~68 (
// Equation(s):
// \rfif.rdat1[28]~68_combout  = (Instr_IF_23 & ((\rfif.rdat1[28]~67_combout  & (\regs[31][28]~q )) # (!\rfif.rdat1[28]~67_combout  & ((\regs[23][28]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[28]~67_combout ))))

	.dataa(\regs[31][28]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[23][28]~q ),
	.datad(\rfif.rdat1[28]~67_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~68_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~68 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[28]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \regs[29][28]~feeder (
// Equation(s):
// \regs[29][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[29][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N7
dffeas \regs[29][28] (
	.clk(!CLK),
	.d(\regs[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][28] .is_wysiwyg = "true";
defparam \regs[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \regs[17][28]~feeder (
// Equation(s):
// \regs[17][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[17][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N27
dffeas \regs[17][28] (
	.clk(!CLK),
	.d(\regs[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][28] .is_wysiwyg = "true";
defparam \regs[17][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N29
dffeas \regs[25][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][28] .is_wysiwyg = "true";
defparam \regs[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[28]~60 (
// Equation(s):
// \rfif.rdat1[28]~60_combout  = (Instr_IF_24 & (((\regs[25][28]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][28]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][28]~q ),
	.datac(\regs[25][28]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~60_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~60 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[28]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N25
dffeas \regs[21][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][28] .is_wysiwyg = "true";
defparam \regs[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[28]~61 (
// Equation(s):
// \rfif.rdat1[28]~61_combout  = (\rfif.rdat1[28]~60_combout  & ((\regs[29][28]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[28]~60_combout  & (((\regs[21][28]~q  & Instr_IF_23))))

	.dataa(\regs[29][28]~q ),
	.datab(\rfif.rdat1[28]~60_combout ),
	.datac(\regs[21][28]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~61_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~61 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[28]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N23
dffeas \regs[15][28] (
	.clk(!CLK),
	.d(input_b2),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][28] .is_wysiwyg = "true";
defparam \regs[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N23
dffeas \regs[14][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][28] .is_wysiwyg = "true";
defparam \regs[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N9
dffeas \regs[13][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][28] .is_wysiwyg = "true";
defparam \regs[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \rfif.rdat1[28]~77 (
// Equation(s):
// \rfif.rdat1[28]~77_combout  = (Instr_IF_21 & (((\regs[13][28]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][28]~q  & ((!Instr_IF_22))))

	.dataa(\regs[12][28]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][28]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~77_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~77 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[28]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \rfif.rdat1[28]~78 (
// Equation(s):
// \rfif.rdat1[28]~78_combout  = (Instr_IF_22 & ((\rfif.rdat1[28]~77_combout  & (\regs[15][28]~q )) # (!\rfif.rdat1[28]~77_combout  & ((\regs[14][28]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[28]~77_combout ))))

	.dataa(\regs[15][28]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[14][28]~q ),
	.datad(\rfif.rdat1[28]~77_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~78_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~78 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[28]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N15
dffeas \regs[9][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][28] .is_wysiwyg = "true";
defparam \regs[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N29
dffeas \regs[11][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][28] .is_wysiwyg = "true";
defparam \regs[11][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[28]~73 (
// Equation(s):
// \rfif.rdat1[28]~73_combout  = (\rfif.rdat1[28]~72_combout  & (((\regs[11][28]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[28]~72_combout  & (Instr_IF_21 & (\regs[9][28]~q )))

	.dataa(\rfif.rdat1[28]~72_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[9][28]~q ),
	.datad(\regs[11][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~73_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~73 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[28]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \regs[2][28]~feeder (
// Equation(s):
// \regs[2][28]~feeder_combout  = \input_b~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][28]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \regs[2][28] (
	.clk(!CLK),
	.d(\regs[2][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][28] .is_wysiwyg = "true";
defparam \regs[2][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N19
dffeas \regs[0][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][28] .is_wysiwyg = "true";
defparam \regs[0][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \rfif.rdat1[28]~74 (
// Equation(s):
// \rfif.rdat1[28]~74_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][28]~q )) # (!Instr_IF_22 & ((\regs[0][28]~q )))))

	.dataa(Instr_IF_21),
	.datab(\regs[2][28]~q ),
	.datac(\regs[0][28]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~74_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~74 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[28]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N7
dffeas \regs[1][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][28] .is_wysiwyg = "true";
defparam \regs[1][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N1
dffeas \regs[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][28] .is_wysiwyg = "true";
defparam \regs[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[28]~75 (
// Equation(s):
// \rfif.rdat1[28]~75_combout  = (Instr_IF_21 & ((\rfif.rdat1[28]~74_combout  & ((\regs[3][28]~q ))) # (!\rfif.rdat1[28]~74_combout  & (\regs[1][28]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[28]~74_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[28]~74_combout ),
	.datac(\regs[1][28]~q ),
	.datad(\regs[3][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~75_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~75 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[28]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \rfif.rdat1[28]~76 (
// Equation(s):
// \rfif.rdat1[28]~76_combout  = (Instr_IF_24 & ((\rfif.rdat1[28]~73_combout ) # ((Instr_IF_23)))) # (!Instr_IF_24 & (((!Instr_IF_23 & \rfif.rdat1[28]~75_combout ))))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[28]~73_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[28]~75_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~76_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~76 .lut_mask = 16'hADA8;
defparam \rfif.rdat1[28]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N3
dffeas \regs[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][28] .is_wysiwyg = "true";
defparam \regs[4][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N27
dffeas \regs[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][28] .is_wysiwyg = "true";
defparam \regs[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[28]~70 (
// Equation(s):
// \rfif.rdat1[28]~70_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][28]~q ))) # (!Instr_IF_21 & (\regs[4][28]~q ))))

	.dataa(Instr_IF_22),
	.datab(\regs[4][28]~q ),
	.datac(\regs[5][28]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~70_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~70 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[28]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N17
dffeas \regs[7][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][28] .is_wysiwyg = "true";
defparam \regs[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N13
dffeas \regs[6][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][28] .is_wysiwyg = "true";
defparam \regs[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[28]~71 (
// Equation(s):
// \rfif.rdat1[28]~71_combout  = (\rfif.rdat1[28]~70_combout  & ((\regs[7][28]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[28]~70_combout  & (((\regs[6][28]~q  & Instr_IF_22))))

	.dataa(\rfif.rdat1[28]~70_combout ),
	.datab(\regs[7][28]~q ),
	.datac(\regs[6][28]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[28]~71_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[28]~71 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[28]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N27
dffeas \regs[12][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][28] .is_wysiwyg = "true";
defparam \regs[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \rfif.rdat2[28]~80 (
// Equation(s):
// \rfif.rdat2[28]~80_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[13][28]~q )) # (!Instr_IF_16 & ((\regs[12][28]~q )))))

	.dataa(\regs[13][28]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[12][28]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~80_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~80 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[28]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[28]~81 (
// Equation(s):
// \rfif.rdat2[28]~81_combout  = (Instr_IF_17 & ((\rfif.rdat2[28]~80_combout  & (\regs[15][28]~q )) # (!\rfif.rdat2[28]~80_combout  & ((\regs[14][28]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[28]~80_combout ))))

	.dataa(\regs[15][28]~q ),
	.datab(\regs[14][28]~q ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[28]~80_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~81_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~81 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[28]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[28]~73 (
// Equation(s):
// \rfif.rdat2[28]~73_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][28]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][28]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][28]~q ),
	.datad(\regs[5][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~73_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~73 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[28]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[28]~74 (
// Equation(s):
// \rfif.rdat2[28]~74_combout  = (Instr_IF_17 & ((\rfif.rdat2[28]~73_combout  & ((\regs[7][28]~q ))) # (!\rfif.rdat2[28]~73_combout  & (\regs[6][28]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[28]~73_combout ))))

	.dataa(\regs[6][28]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[7][28]~q ),
	.datad(\rfif.rdat2[28]~73_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~74_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~74 .lut_mask = 16'hF388;
defparam \rfif.rdat2[28]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \rfif.rdat2[28]~77 (
// Equation(s):
// \rfif.rdat2[28]~77_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][28]~q )) # (!Instr_IF_17 & ((\regs[0][28]~q )))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[2][28]~q ),
	.datad(\regs[0][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~77_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~77 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[28]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \rfif.rdat2[28]~78 (
// Equation(s):
// \rfif.rdat2[28]~78_combout  = (Instr_IF_16 & ((\rfif.rdat2[28]~77_combout  & (\regs[3][28]~q )) # (!\rfif.rdat2[28]~77_combout  & ((\regs[1][28]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[28]~77_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[28]~77_combout ),
	.datac(\regs[3][28]~q ),
	.datad(\regs[1][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~78_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~78 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[28]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N23
dffeas \regs[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][28] .is_wysiwyg = "true";
defparam \regs[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N29
dffeas \regs[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][28] .is_wysiwyg = "true";
defparam \regs[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[28]~75 (
// Equation(s):
// \rfif.rdat2[28]~75_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][28]~q ))) # (!Instr_IF_17 & (\regs[8][28]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][28]~q ),
	.datad(\regs[10][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~75_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~75 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[28]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[28]~76 (
// Equation(s):
// \rfif.rdat2[28]~76_combout  = (Instr_IF_16 & ((\rfif.rdat2[28]~75_combout  & ((\regs[11][28]~q ))) # (!\rfif.rdat2[28]~75_combout  & (\regs[9][28]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[28]~75_combout ))))

	.dataa(\regs[9][28]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[11][28]~q ),
	.datad(\rfif.rdat2[28]~75_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~76_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~76 .lut_mask = 16'hF388;
defparam \rfif.rdat2[28]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[28]~79 (
// Equation(s):
// \rfif.rdat2[28]~79_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\rfif.rdat2[28]~76_combout )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\rfif.rdat2[28]~78_combout )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[28]~78_combout ),
	.datad(\rfif.rdat2[28]~76_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~79_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~79 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[28]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \rfif.rdat2[28]~82 (
// Equation(s):
// \rfif.rdat2[28]~82_combout  = (Instr_IF_18 & ((\rfif.rdat2[28]~79_combout  & (\rfif.rdat2[28]~81_combout )) # (!\rfif.rdat2[28]~79_combout  & ((\rfif.rdat2[28]~74_combout ))))) # (!Instr_IF_18 & (((\rfif.rdat2[28]~79_combout ))))

	.dataa(\rfif.rdat2[28]~81_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[28]~74_combout ),
	.datad(\rfif.rdat2[28]~79_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~82_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~82 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[28]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \rfif.rdat2[28]~70 (
// Equation(s):
// \rfif.rdat2[28]~70_combout  = (Instr_IF_19 & ((\regs[27][28]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[19][28]~q  & !Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][28]~q ),
	.datac(\regs[19][28]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~70_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~70 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[28]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \rfif.rdat2[28]~71 (
// Equation(s):
// \rfif.rdat2[28]~71_combout  = (Instr_IF_18 & ((\rfif.rdat2[28]~70_combout  & (\regs[31][28]~q )) # (!\rfif.rdat2[28]~70_combout  & ((\regs[23][28]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[28]~70_combout ))))

	.dataa(\regs[31][28]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[23][28]~q ),
	.datad(\rfif.rdat2[28]~70_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~71_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~71 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[28]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \rfif.rdat2[28]~63 (
// Equation(s):
// \rfif.rdat2[28]~63_combout  = (Instr_IF_19 & (((Instr_IF_18) # (\regs[25][28]~q )))) # (!Instr_IF_19 & (\regs[17][28]~q  & (!Instr_IF_18)))

	.dataa(Instr_IF_19),
	.datab(\regs[17][28]~q ),
	.datac(Instr_IF_18),
	.datad(\regs[25][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~63_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~63 .lut_mask = 16'hAEA4;
defparam \rfif.rdat2[28]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[28]~64 (
// Equation(s):
// \rfif.rdat2[28]~64_combout  = (\rfif.rdat2[28]~63_combout  & ((\regs[29][28]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[28]~63_combout  & (((Instr_IF_18 & \regs[21][28]~q ))))

	.dataa(\regs[29][28]~q ),
	.datab(\rfif.rdat2[28]~63_combout ),
	.datac(Instr_IF_18),
	.datad(\regs[21][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~64_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~64 .lut_mask = 16'hBC8C;
defparam \rfif.rdat2[28]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[28]~67 (
// Equation(s):
// \rfif.rdat2[28]~67_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][28]~q ))) # (!Instr_IF_18 & (\regs[16][28]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][28]~q ),
	.datad(\regs[20][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~67_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~67 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[28]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[28]~68 (
// Equation(s):
// \rfif.rdat2[28]~68_combout  = (Instr_IF_19 & ((\rfif.rdat2[28]~67_combout  & (\regs[28][28]~q )) # (!\rfif.rdat2[28]~67_combout  & ((\regs[24][28]~q ))))) # (!Instr_IF_19 & (((\rfif.rdat2[28]~67_combout ))))

	.dataa(\regs[28][28]~q ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[28]~67_combout ),
	.datad(\regs[24][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~68_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~68 .lut_mask = 16'hBCB0;
defparam \rfif.rdat2[28]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \regs[18][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][28] .is_wysiwyg = "true";
defparam \regs[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \rfif.rdat2[28]~65 (
// Equation(s):
// \rfif.rdat2[28]~65_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][28]~q ))) # (!Instr_IF_18 & (\regs[18][28]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][28]~q ),
	.datad(\regs[22][28]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~65_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~65 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[28]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[28]~66 (
// Equation(s):
// \rfif.rdat2[28]~66_combout  = (Instr_IF_19 & ((\rfif.rdat2[28]~65_combout  & ((\regs[30][28]~q ))) # (!\rfif.rdat2[28]~65_combout  & (\regs[26][28]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[28]~65_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][28]~q ),
	.datac(\regs[30][28]~q ),
	.datad(\rfif.rdat2[28]~65_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~66_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~66 .lut_mask = 16'hF588;
defparam \rfif.rdat2[28]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[28]~69 (
// Equation(s):
// \rfif.rdat2[28]~69_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[28]~66_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[28]~68_combout ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[28]~68_combout ),
	.datad(\rfif.rdat2[28]~66_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~69_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~69 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[28]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[28]~72 (
// Equation(s):
// \rfif.rdat2[28]~72_combout  = (Instr_IF_16 & ((\rfif.rdat2[28]~69_combout  & (\rfif.rdat2[28]~71_combout )) # (!\rfif.rdat2[28]~69_combout  & ((\rfif.rdat2[28]~64_combout ))))) # (!Instr_IF_16 & (((\rfif.rdat2[28]~69_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[28]~71_combout ),
	.datac(\rfif.rdat2[28]~64_combout ),
	.datad(\rfif.rdat2[28]~69_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[28]~72_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[28]~72 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[28]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \regs[23][27]~feeder (
// Equation(s):
// \regs[23][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b3),
	.cin(gnd),
	.combout(\regs[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][27]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N19
dffeas \regs[23][27] (
	.clk(!CLK),
	.d(\regs[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][27] .is_wysiwyg = "true";
defparam \regs[23][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N7
dffeas \regs[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][27] .is_wysiwyg = "true";
defparam \regs[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[27]~87 (
// Equation(s):
// \rfif.rdat1[27]~87_combout  = (Instr_IF_23 & ((\regs[23][27]~q ) # ((Instr_IF_24)))) # (!Instr_IF_23 & (((!Instr_IF_24 & \regs[19][27]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[23][27]~q ),
	.datac(Instr_IF_24),
	.datad(\regs[19][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~87_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~87 .lut_mask = 16'hADA8;
defparam \rfif.rdat1[27]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N25
dffeas \regs[31][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][27] .is_wysiwyg = "true";
defparam \regs[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N3
dffeas \regs[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][27] .is_wysiwyg = "true";
defparam \regs[27][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[27]~88 (
// Equation(s):
// \rfif.rdat1[27]~88_combout  = (\rfif.rdat1[27]~87_combout  & ((\regs[31][27]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[27]~87_combout  & (((\regs[27][27]~q  & Instr_IF_24))))

	.dataa(\rfif.rdat1[27]~87_combout ),
	.datab(\regs[31][27]~q ),
	.datac(\regs[27][27]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~88_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~88 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[27]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N9
dffeas \regs[22][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][27] .is_wysiwyg = "true";
defparam \regs[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \regs[30][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][27] .is_wysiwyg = "true";
defparam \regs[30][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \regs[18][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][27] .is_wysiwyg = "true";
defparam \regs[18][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N3
dffeas \regs[26][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][27] .is_wysiwyg = "true";
defparam \regs[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \rfif.rdat1[27]~80 (
// Equation(s):
// \rfif.rdat1[27]~80_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[26][27]~q ))) # (!Instr_IF_24 & (\regs[18][27]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[18][27]~q ),
	.datac(\regs[26][27]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~80_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~80 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[27]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \rfif.rdat1[27]~81 (
// Equation(s):
// \rfif.rdat1[27]~81_combout  = (Instr_IF_23 & ((\rfif.rdat1[27]~80_combout  & ((\regs[30][27]~q ))) # (!\rfif.rdat1[27]~80_combout  & (\regs[22][27]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[27]~80_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[22][27]~q ),
	.datac(\regs[30][27]~q ),
	.datad(\rfif.rdat1[27]~80_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~81_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~81 .lut_mask = 16'hF588;
defparam \rfif.rdat1[27]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N20
cycloneive_lcell_comb \regs[20][27]~feeder (
// Equation(s):
// \regs[20][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b3),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N21
dffeas \regs[20][27] (
	.clk(!CLK),
	.d(\regs[20][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][27] .is_wysiwyg = "true";
defparam \regs[20][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N9
dffeas \regs[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][27] .is_wysiwyg = "true";
defparam \regs[16][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N19
dffeas \regs[24][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][27] .is_wysiwyg = "true";
defparam \regs[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[27]~84 (
// Equation(s):
// \rfif.rdat1[27]~84_combout  = (Instr_IF_24 & (((\regs[24][27]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[16][27]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[16][27]~q ),
	.datac(\regs[24][27]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~84_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~84 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[27]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[27]~85 (
// Equation(s):
// \rfif.rdat1[27]~85_combout  = (\rfif.rdat1[27]~84_combout  & ((\regs[28][27]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[27]~84_combout  & (((\regs[20][27]~q  & Instr_IF_23))))

	.dataa(\regs[28][27]~q ),
	.datab(\regs[20][27]~q ),
	.datac(\rfif.rdat1[27]~84_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~85_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~85 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[27]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \regs[25][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][27] .is_wysiwyg = "true";
defparam \regs[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N15
dffeas \regs[17][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][27] .is_wysiwyg = "true";
defparam \regs[17][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N17
dffeas \regs[21][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][27] .is_wysiwyg = "true";
defparam \regs[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[27]~82 (
// Equation(s):
// \rfif.rdat1[27]~82_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][27]~q ))) # (!Instr_IF_23 & (\regs[17][27]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][27]~q ),
	.datac(\regs[21][27]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~82_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~82 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[27]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[27]~83 (
// Equation(s):
// \rfif.rdat1[27]~83_combout  = (Instr_IF_24 & ((\rfif.rdat1[27]~82_combout  & (\regs[29][27]~q )) # (!\rfif.rdat1[27]~82_combout  & ((\regs[25][27]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[27]~82_combout ))))

	.dataa(\regs[29][27]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[25][27]~q ),
	.datad(\rfif.rdat1[27]~82_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~83_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~83 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[27]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[27]~86 (
// Equation(s):
// \rfif.rdat1[27]~86_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & ((\rfif.rdat1[27]~83_combout ))) # (!Instr_IF_21 & (\rfif.rdat1[27]~85_combout ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[27]~85_combout ),
	.datad(\rfif.rdat1[27]~83_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~86_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~86 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[27]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \regs[1][27]~feeder (
// Equation(s):
// \regs[1][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b3),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[1][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[1][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N1
dffeas \regs[1][27] (
	.clk(!CLK),
	.d(\regs[1][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][27] .is_wysiwyg = "true";
defparam \regs[1][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N17
dffeas \regs[0][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][27] .is_wysiwyg = "true";
defparam \regs[0][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[27]~94 (
// Equation(s):
// \rfif.rdat1[27]~94_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][27]~q )) # (!Instr_IF_21 & ((\regs[0][27]~q )))))

	.dataa(Instr_IF_22),
	.datab(\regs[1][27]~q ),
	.datac(\regs[0][27]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~94_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~94 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[27]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N23
dffeas \regs[2][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][27] .is_wysiwyg = "true";
defparam \regs[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N13
dffeas \regs[3][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][27] .is_wysiwyg = "true";
defparam \regs[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \rfif.rdat1[27]~95 (
// Equation(s):
// \rfif.rdat1[27]~95_combout  = (Instr_IF_22 & ((\rfif.rdat1[27]~94_combout  & ((\regs[3][27]~q ))) # (!\rfif.rdat1[27]~94_combout  & (\regs[2][27]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[27]~94_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[27]~94_combout ),
	.datac(\regs[2][27]~q ),
	.datad(\regs[3][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~95_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~95 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[27]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N13
dffeas \regs[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][27] .is_wysiwyg = "true";
defparam \regs[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N7
dffeas \regs[7][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][27] .is_wysiwyg = "true";
defparam \regs[7][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[27]~93 (
// Equation(s):
// \rfif.rdat1[27]~93_combout  = (\rfif.rdat1[27]~92_combout  & (((\regs[7][27]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[27]~92_combout  & (Instr_IF_21 & (\regs[5][27]~q )))

	.dataa(\rfif.rdat1[27]~92_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[5][27]~q ),
	.datad(\regs[7][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~93_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~93 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[27]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[27]~96 (
// Equation(s):
// \rfif.rdat1[27]~96_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\rfif.rdat1[27]~93_combout ))) # (!Instr_IF_23 & (\rfif.rdat1[27]~95_combout ))))

	.dataa(\rfif.rdat1[27]~95_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[27]~93_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~96_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~96 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[27]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \regs[15][27]~feeder (
// Equation(s):
// \regs[15][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b3),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N5
dffeas \regs[15][27] (
	.clk(!CLK),
	.d(\regs[15][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][27] .is_wysiwyg = "true";
defparam \regs[15][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N9
dffeas \regs[13][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][27] .is_wysiwyg = "true";
defparam \regs[13][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \regs[14][27]~feeder (
// Equation(s):
// \regs[14][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b3),
	.cin(gnd),
	.combout(\regs[14][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][27]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N5
dffeas \regs[14][27] (
	.clk(!CLK),
	.d(\regs[14][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][27] .is_wysiwyg = "true";
defparam \regs[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N15
dffeas \regs[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][27] .is_wysiwyg = "true";
defparam \regs[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[27]~97 (
// Equation(s):
// \rfif.rdat1[27]~97_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[14][27]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[12][27]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[14][27]~q ),
	.datad(\regs[12][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~97_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~97 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[27]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[27]~98 (
// Equation(s):
// \rfif.rdat1[27]~98_combout  = (Instr_IF_21 & ((\rfif.rdat1[27]~97_combout  & (\regs[15][27]~q )) # (!\rfif.rdat1[27]~97_combout  & ((\regs[13][27]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[27]~97_combout ))))

	.dataa(\regs[15][27]~q ),
	.datab(\regs[13][27]~q ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[27]~97_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~98_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~98 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[27]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \regs[11][27]~feeder (
// Equation(s):
// \regs[11][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b3),
	.cin(gnd),
	.combout(\regs[11][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][27]~feeder .lut_mask = 16'hFF00;
defparam \regs[11][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N5
dffeas \regs[11][27] (
	.clk(!CLK),
	.d(\regs[11][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][27] .is_wysiwyg = "true";
defparam \regs[11][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \regs[10][27]~feeder (
// Equation(s):
// \regs[10][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b3),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N19
dffeas \regs[10][27] (
	.clk(!CLK),
	.d(\regs[10][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][27] .is_wysiwyg = "true";
defparam \regs[10][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N23
dffeas \regs[9][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][27] .is_wysiwyg = "true";
defparam \regs[9][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N29
dffeas \regs[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][27] .is_wysiwyg = "true";
defparam \regs[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N22
cycloneive_lcell_comb \rfif.rdat1[27]~90 (
// Equation(s):
// \rfif.rdat1[27]~90_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][27]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[8][27]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[9][27]~q ),
	.datad(\regs[8][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~90_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~90 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[27]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[27]~91 (
// Equation(s):
// \rfif.rdat1[27]~91_combout  = (Instr_IF_22 & ((\rfif.rdat1[27]~90_combout  & (\regs[11][27]~q )) # (!\rfif.rdat1[27]~90_combout  & ((\regs[10][27]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[27]~90_combout ))))

	.dataa(\regs[11][27]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[10][27]~q ),
	.datad(\rfif.rdat1[27]~90_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[27]~91_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[27]~91 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[27]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[27]~94 (
// Equation(s):
// \rfif.rdat2[27]~94_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][27]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][27]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][27]~q ),
	.datad(\regs[9][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~94_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~94 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[27]~95 (
// Equation(s):
// \rfif.rdat2[27]~95_combout  = (\rfif.rdat2[27]~94_combout  & ((\regs[11][27]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[27]~94_combout  & (((Instr_IF_17 & \regs[10][27]~q ))))

	.dataa(\regs[11][27]~q ),
	.datab(\rfif.rdat2[27]~94_combout ),
	.datac(Instr_IF_17),
	.datad(\regs[10][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~95_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~95 .lut_mask = 16'hBC8C;
defparam \rfif.rdat2[27]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[27]~101 (
// Equation(s):
// \rfif.rdat2[27]~101_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][27]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][27]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][27]~q ),
	.datad(\regs[14][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~101_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~101 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[27]~102 (
// Equation(s):
// \rfif.rdat2[27]~102_combout  = (\rfif.rdat2[27]~101_combout  & ((\regs[15][27]~q ) # ((!Instr_IF_16)))) # (!\rfif.rdat2[27]~101_combout  & (((\regs[13][27]~q  & Instr_IF_16))))

	.dataa(\regs[15][27]~q ),
	.datab(\rfif.rdat2[27]~101_combout ),
	.datac(\regs[13][27]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~102_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~102 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[27]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N13
dffeas \regs[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][27] .is_wysiwyg = "true";
defparam \regs[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[27]~96 (
// Equation(s):
// \rfif.rdat2[27]~96_combout  = (Instr_IF_17 & ((\regs[6][27]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\regs[4][27]~q  & !Instr_IF_16))))

	.dataa(\regs[6][27]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[4][27]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~96_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~96 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[27]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[27]~97 (
// Equation(s):
// \rfif.rdat2[27]~97_combout  = (Instr_IF_16 & ((\rfif.rdat2[27]~96_combout  & (\regs[7][27]~q )) # (!\rfif.rdat2[27]~96_combout  & ((\regs[5][27]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[27]~96_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[27]~96_combout ),
	.datac(\regs[7][27]~q ),
	.datad(\regs[5][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~97_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~97 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[27]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \rfif.rdat2[27]~98 (
// Equation(s):
// \rfif.rdat2[27]~98_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[1][27]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[0][27]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][27]~q ),
	.datad(\regs[1][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~98_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~98 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \rfif.rdat2[27]~99 (
// Equation(s):
// \rfif.rdat2[27]~99_combout  = (Instr_IF_17 & ((\rfif.rdat2[27]~98_combout  & ((\regs[3][27]~q ))) # (!\rfif.rdat2[27]~98_combout  & (\regs[2][27]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[27]~98_combout ))))

	.dataa(\regs[2][27]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[3][27]~q ),
	.datad(\rfif.rdat2[27]~98_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~99_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~99 .lut_mask = 16'hF388;
defparam \rfif.rdat2[27]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[27]~100 (
// Equation(s):
// \rfif.rdat2[27]~100_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\rfif.rdat2[27]~97_combout )))) # (!Instr_IF_18 & (!Instr_IF_19 & ((\rfif.rdat2[27]~99_combout ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[27]~97_combout ),
	.datad(\rfif.rdat2[27]~99_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~100_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~100 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[27]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \rfif.rdat2[27]~103 (
// Equation(s):
// \rfif.rdat2[27]~103_combout  = (\rfif.rdat2[27]~100_combout  & (((\rfif.rdat2[27]~102_combout ) # (!Instr_IF_19)))) # (!\rfif.rdat2[27]~100_combout  & (\rfif.rdat2[27]~95_combout  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[27]~95_combout ),
	.datab(\rfif.rdat2[27]~102_combout ),
	.datac(\rfif.rdat2[27]~100_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~103_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~103 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[27]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[27]~91 (
// Equation(s):
// \rfif.rdat2[27]~91_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[23][27]~q )) # (!Instr_IF_18 & ((\regs[19][27]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[23][27]~q ),
	.datac(\regs[19][27]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~91_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~91 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[27]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N24
cycloneive_lcell_comb \rfif.rdat2[27]~92 (
// Equation(s):
// \rfif.rdat2[27]~92_combout  = (Instr_IF_19 & ((\rfif.rdat2[27]~91_combout  & ((\regs[31][27]~q ))) # (!\rfif.rdat2[27]~91_combout  & (\regs[27][27]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[27]~91_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][27]~q ),
	.datac(\regs[31][27]~q ),
	.datad(\rfif.rdat2[27]~91_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~92_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~92 .lut_mask = 16'hF588;
defparam \rfif.rdat2[27]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[27]~84 (
// Equation(s):
// \rfif.rdat2[27]~84_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][27]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][27]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][27]~q ),
	.datad(\regs[26][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~84_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~84 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \rfif.rdat2[27]~85 (
// Equation(s):
// \rfif.rdat2[27]~85_combout  = (\rfif.rdat2[27]~84_combout  & ((\regs[30][27]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[27]~84_combout  & (((\regs[22][27]~q  & Instr_IF_18))))

	.dataa(\regs[30][27]~q ),
	.datab(\rfif.rdat2[27]~84_combout ),
	.datac(\regs[22][27]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~85_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~85 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[27]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \regs[29][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][27] .is_wysiwyg = "true";
defparam \regs[29][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[27]~86 (
// Equation(s):
// \rfif.rdat2[27]~86_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[21][27]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[17][27]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][27]~q ),
	.datad(\regs[21][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~86_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~86 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[27]~87 (
// Equation(s):
// \rfif.rdat2[27]~87_combout  = (Instr_IF_19 & ((\rfif.rdat2[27]~86_combout  & ((\regs[29][27]~q ))) # (!\rfif.rdat2[27]~86_combout  & (\regs[25][27]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[27]~86_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][27]~q ),
	.datac(\regs[29][27]~q ),
	.datad(\rfif.rdat2[27]~86_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~87_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~87 .lut_mask = 16'hF588;
defparam \rfif.rdat2[27]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N14
cycloneive_lcell_comb \regs[28][27]~feeder (
// Equation(s):
// \regs[28][27]~feeder_combout  = \input_b~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b3),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][27]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N15
dffeas \regs[28][27] (
	.clk(!CLK),
	.d(\regs[28][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][27] .is_wysiwyg = "true";
defparam \regs[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[27]~88 (
// Equation(s):
// \rfif.rdat2[27]~88_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[24][27]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[16][27]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][27]~q ),
	.datad(\regs[24][27]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~88_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~88 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[27]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[27]~89 (
// Equation(s):
// \rfif.rdat2[27]~89_combout  = (Instr_IF_18 & ((\rfif.rdat2[27]~88_combout  & ((\regs[28][27]~q ))) # (!\rfif.rdat2[27]~88_combout  & (\regs[20][27]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[27]~88_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[20][27]~q ),
	.datac(\regs[28][27]~q ),
	.datad(\rfif.rdat2[27]~88_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~89_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~89 .lut_mask = 16'hF588;
defparam \rfif.rdat2[27]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[27]~90 (
// Equation(s):
// \rfif.rdat2[27]~90_combout  = (Instr_IF_16 & ((\rfif.rdat2[27]~87_combout ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((!Instr_IF_17 & \rfif.rdat2[27]~89_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[27]~87_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[27]~89_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~90_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~90 .lut_mask = 16'hADA8;
defparam \rfif.rdat2[27]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \rfif.rdat2[27]~93 (
// Equation(s):
// \rfif.rdat2[27]~93_combout  = (Instr_IF_17 & ((\rfif.rdat2[27]~90_combout  & (\rfif.rdat2[27]~92_combout )) # (!\rfif.rdat2[27]~90_combout  & ((\rfif.rdat2[27]~85_combout ))))) # (!Instr_IF_17 & (((\rfif.rdat2[27]~90_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[27]~92_combout ),
	.datac(\rfif.rdat2[27]~85_combout ),
	.datad(\rfif.rdat2[27]~90_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[27]~93_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[27]~93 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[27]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N27
dffeas \regs[31][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][26] .is_wysiwyg = "true";
defparam \regs[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \regs[23][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][26] .is_wysiwyg = "true";
defparam \regs[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N3
dffeas \regs[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][26] .is_wysiwyg = "true";
defparam \regs[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \regs[27][26]~feeder (
// Equation(s):
// \regs[27][26]~feeder_combout  = \input_b~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b4),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][26]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N5
dffeas \regs[27][26] (
	.clk(!CLK),
	.d(\regs[27][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][26] .is_wysiwyg = "true";
defparam \regs[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[26]~107 (
// Equation(s):
// \rfif.rdat1[26]~107_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[27][26]~q ))) # (!Instr_IF_24 & (\regs[19][26]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[19][26]~q ),
	.datad(\regs[27][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~107_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~107 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[26]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[26]~108 (
// Equation(s):
// \rfif.rdat1[26]~108_combout  = (Instr_IF_23 & ((\rfif.rdat1[26]~107_combout  & (\regs[31][26]~q )) # (!\rfif.rdat1[26]~107_combout  & ((\regs[23][26]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[26]~107_combout ))))

	.dataa(\regs[31][26]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[23][26]~q ),
	.datad(\rfif.rdat1[26]~107_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~108_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~108 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[26]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N9
dffeas \regs[21][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][26] .is_wysiwyg = "true";
defparam \regs[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N27
dffeas \regs[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][26] .is_wysiwyg = "true";
defparam \regs[17][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N9
dffeas \regs[25][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][26] .is_wysiwyg = "true";
defparam \regs[25][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \rfif.rdat1[26]~100 (
// Equation(s):
// \rfif.rdat1[26]~100_combout  = (Instr_IF_24 & (((\regs[25][26]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][26]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][26]~q ),
	.datac(\regs[25][26]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~100_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~100 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[26]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N31
dffeas \regs[29][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][26] .is_wysiwyg = "true";
defparam \regs[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \rfif.rdat1[26]~101 (
// Equation(s):
// \rfif.rdat1[26]~101_combout  = (\rfif.rdat1[26]~100_combout  & (((\regs[29][26]~q ) # (!Instr_IF_23)))) # (!\rfif.rdat1[26]~100_combout  & (\regs[21][26]~q  & ((Instr_IF_23))))

	.dataa(\regs[21][26]~q ),
	.datab(\rfif.rdat1[26]~100_combout ),
	.datac(\regs[29][26]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~101_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~101 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[26]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N21
dffeas \regs[16][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][26] .is_wysiwyg = "true";
defparam \regs[16][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N3
dffeas \regs[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][26] .is_wysiwyg = "true";
defparam \regs[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[26]~104 (
// Equation(s):
// \rfif.rdat1[26]~104_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[20][26]~q ))) # (!Instr_IF_23 & (\regs[16][26]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[16][26]~q ),
	.datac(\regs[20][26]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~104_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~104 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[26]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y39_N3
dffeas \regs[24][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][26] .is_wysiwyg = "true";
defparam \regs[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N21
dffeas \regs[28][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][26] .is_wysiwyg = "true";
defparam \regs[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[26]~105 (
// Equation(s):
// \rfif.rdat1[26]~105_combout  = (Instr_IF_24 & ((\rfif.rdat1[26]~104_combout  & ((\regs[28][26]~q ))) # (!\rfif.rdat1[26]~104_combout  & (\regs[24][26]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[26]~104_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[26]~104_combout ),
	.datac(\regs[24][26]~q ),
	.datad(\regs[28][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~105_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~105 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[26]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N19
dffeas \regs[30][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][26] .is_wysiwyg = "true";
defparam \regs[30][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N9
dffeas \regs[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][26] .is_wysiwyg = "true";
defparam \regs[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N1
dffeas \regs[22][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][26] .is_wysiwyg = "true";
defparam \regs[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[26]~102 (
// Equation(s):
// \rfif.rdat1[26]~102_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][26]~q ))) # (!Instr_IF_23 & (\regs[18][26]~q ))))

	.dataa(\regs[18][26]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[22][26]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~102_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~102 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[26]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[26]~103 (
// Equation(s):
// \rfif.rdat1[26]~103_combout  = (Instr_IF_24 & ((\rfif.rdat1[26]~102_combout  & (\regs[30][26]~q )) # (!\rfif.rdat1[26]~102_combout  & ((\regs[26][26]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[26]~102_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[30][26]~q ),
	.datac(\regs[26][26]~q ),
	.datad(\rfif.rdat1[26]~102_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~103_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~103 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[26]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \rfif.rdat1[26]~106 (
// Equation(s):
// \rfif.rdat1[26]~106_combout  = (Instr_IF_22 & (((\rfif.rdat1[26]~103_combout ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\rfif.rdat1[26]~105_combout  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[26]~105_combout ),
	.datac(\rfif.rdat1[26]~103_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~106_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~106 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[26]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N25
dffeas \regs[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][26] .is_wysiwyg = "true";
defparam \regs[6][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N21
dffeas \regs[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][26] .is_wysiwyg = "true";
defparam \regs[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N3
dffeas \regs[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][26] .is_wysiwyg = "true";
defparam \regs[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[26]~110 (
// Equation(s):
// \rfif.rdat1[26]~110_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][26]~q ))) # (!Instr_IF_21 & (\regs[4][26]~q ))))

	.dataa(\regs[4][26]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][26]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~110_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~110 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[26]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[26]~111 (
// Equation(s):
// \rfif.rdat1[26]~111_combout  = (Instr_IF_22 & ((\rfif.rdat1[26]~110_combout  & ((\regs[7][26]~q ))) # (!\rfif.rdat1[26]~110_combout  & (\regs[6][26]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[26]~110_combout ))))

	.dataa(\regs[6][26]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[7][26]~q ),
	.datad(\rfif.rdat1[26]~110_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~111_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~111 .lut_mask = 16'hF388;
defparam \rfif.rdat1[26]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \regs[14][26]~feeder (
// Equation(s):
// \regs[14][26]~feeder_combout  = \input_b~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b4),
	.cin(gnd),
	.combout(\regs[14][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][26]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N3
dffeas \regs[14][26] (
	.clk(!CLK),
	.d(\regs[14][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][26] .is_wysiwyg = "true";
defparam \regs[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N23
dffeas \regs[15][26] (
	.clk(!CLK),
	.d(input_b4),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][26] .is_wysiwyg = "true";
defparam \regs[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N15
dffeas \regs[12][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][26] .is_wysiwyg = "true";
defparam \regs[12][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \regs[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][26] .is_wysiwyg = "true";
defparam \regs[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \rfif.rdat1[26]~117 (
// Equation(s):
// \rfif.rdat1[26]~117_combout  = (Instr_IF_21 & (((\regs[13][26]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][26]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][26]~q ),
	.datac(\regs[13][26]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~117_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~117 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[26]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[26]~118 (
// Equation(s):
// \rfif.rdat1[26]~118_combout  = (Instr_IF_22 & ((\rfif.rdat1[26]~117_combout  & ((\regs[15][26]~q ))) # (!\rfif.rdat1[26]~117_combout  & (\regs[14][26]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[26]~117_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[14][26]~q ),
	.datac(\regs[15][26]~q ),
	.datad(\rfif.rdat1[26]~117_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~118_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~118 .lut_mask = 16'hF588;
defparam \rfif.rdat1[26]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N1
dffeas \regs[0][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][26] .is_wysiwyg = "true";
defparam \regs[0][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N31
dffeas \regs[2][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][26] .is_wysiwyg = "true";
defparam \regs[2][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \rfif.rdat1[26]~114 (
// Equation(s):
// \rfif.rdat1[26]~114_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[2][26]~q ))) # (!Instr_IF_22 & (\regs[0][26]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[0][26]~q ),
	.datac(\regs[2][26]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~114_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~114 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[26]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \regs[1][26]~feeder (
// Equation(s):
// \regs[1][26]~feeder_combout  = \input_b~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b4),
	.cin(gnd),
	.combout(\regs[1][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][26]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N25
dffeas \regs[1][26] (
	.clk(!CLK),
	.d(\regs[1][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][26] .is_wysiwyg = "true";
defparam \regs[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[26]~115 (
// Equation(s):
// \rfif.rdat1[26]~115_combout  = (\rfif.rdat1[26]~114_combout  & ((\regs[3][26]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[26]~114_combout  & (((Instr_IF_21 & \regs[1][26]~q ))))

	.dataa(\regs[3][26]~q ),
	.datab(\rfif.rdat1[26]~114_combout ),
	.datac(Instr_IF_21),
	.datad(\regs[1][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~115_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~115 .lut_mask = 16'hBC8C;
defparam \rfif.rdat1[26]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N9
dffeas \regs[11][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][26] .is_wysiwyg = "true";
defparam \regs[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N25
dffeas \regs[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][26] .is_wysiwyg = "true";
defparam \regs[10][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N31
dffeas \regs[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][26] .is_wysiwyg = "true";
defparam \regs[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[26]~112 (
// Equation(s):
// \rfif.rdat1[26]~112_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][26]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][26]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][26]~q ),
	.datad(\regs[8][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~112_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~112 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[26]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N2
cycloneive_lcell_comb \regs[9][26]~feeder (
// Equation(s):
// \regs[9][26]~feeder_combout  = \input_b~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b4),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][26]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N3
dffeas \regs[9][26] (
	.clk(!CLK),
	.d(\regs[9][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][26] .is_wysiwyg = "true";
defparam \regs[9][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \rfif.rdat1[26]~113 (
// Equation(s):
// \rfif.rdat1[26]~113_combout  = (Instr_IF_21 & ((\rfif.rdat1[26]~112_combout  & (\regs[11][26]~q )) # (!\rfif.rdat1[26]~112_combout  & ((\regs[9][26]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[26]~112_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][26]~q ),
	.datac(\rfif.rdat1[26]~112_combout ),
	.datad(\regs[9][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~113_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~113 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[26]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[26]~116 (
// Equation(s):
// \rfif.rdat1[26]~116_combout  = (Instr_IF_24 & (((Instr_IF_23) # (\rfif.rdat1[26]~113_combout )))) # (!Instr_IF_24 & (\rfif.rdat1[26]~115_combout  & (!Instr_IF_23)))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[26]~115_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[26]~113_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[26]~116_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[26]~116 .lut_mask = 16'hAEA4;
defparam \rfif.rdat1[26]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N11
dffeas \regs[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][26] .is_wysiwyg = "true";
defparam \regs[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[26]~115 (
// Equation(s):
// \rfif.rdat2[26]~115_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][26]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][26]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][26]~q ),
	.datad(\regs[5][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~115_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~115 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[26]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \rfif.rdat2[26]~116 (
// Equation(s):
// \rfif.rdat2[26]~116_combout  = (Instr_IF_17 & ((\rfif.rdat2[26]~115_combout  & (\regs[7][26]~q )) # (!\rfif.rdat2[26]~115_combout  & ((\regs[6][26]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[26]~115_combout ))))

	.dataa(\regs[7][26]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[6][26]~q ),
	.datad(\rfif.rdat2[26]~115_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~116_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~116 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[26]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \rfif.rdat2[26]~123 (
// Equation(s):
// \rfif.rdat2[26]~123_combout  = (\rfif.rdat2[26]~122_combout  & (((\regs[15][26]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[26]~122_combout  & (\regs[14][26]~q  & ((Instr_IF_17))))

	.dataa(\rfif.rdat2[26]~122_combout ),
	.datab(\regs[14][26]~q ),
	.datac(\regs[15][26]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~123_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~123 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[26]~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[26]~117 (
// Equation(s):
// \rfif.rdat2[26]~117_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][26]~q ))) # (!Instr_IF_17 & (\regs[8][26]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][26]~q ),
	.datad(\regs[10][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~117_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~117 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[26]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \rfif.rdat2[26]~118 (
// Equation(s):
// \rfif.rdat2[26]~118_combout  = (Instr_IF_16 & ((\rfif.rdat2[26]~117_combout  & ((\regs[11][26]~q ))) # (!\rfif.rdat2[26]~117_combout  & (\regs[9][26]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[26]~117_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][26]~q ),
	.datac(\regs[11][26]~q ),
	.datad(\rfif.rdat2[26]~117_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~118_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~118 .lut_mask = 16'hF588;
defparam \rfif.rdat2[26]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \rfif.rdat2[26]~119 (
// Equation(s):
// \rfif.rdat2[26]~119_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][26]~q )) # (!Instr_IF_17 & ((\regs[0][26]~q )))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[2][26]~q ),
	.datad(\regs[0][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~119_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~119 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[26]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[26]~120 (
// Equation(s):
// \rfif.rdat2[26]~120_combout  = (\rfif.rdat2[26]~119_combout  & ((\regs[3][26]~q ) # ((!Instr_IF_16)))) # (!\rfif.rdat2[26]~119_combout  & (((\regs[1][26]~q  & Instr_IF_16))))

	.dataa(\regs[3][26]~q ),
	.datab(\regs[1][26]~q ),
	.datac(\rfif.rdat2[26]~119_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~120_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~120 .lut_mask = 16'hACF0;
defparam \rfif.rdat2[26]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \rfif.rdat2[26]~121 (
// Equation(s):
// \rfif.rdat2[26]~121_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[26]~118_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[26]~120_combout )))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[26]~118_combout ),
	.datad(\rfif.rdat2[26]~120_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~121_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~121 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[26]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \rfif.rdat2[26]~124 (
// Equation(s):
// \rfif.rdat2[26]~124_combout  = (Instr_IF_18 & ((\rfif.rdat2[26]~121_combout  & ((\rfif.rdat2[26]~123_combout ))) # (!\rfif.rdat2[26]~121_combout  & (\rfif.rdat2[26]~116_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[26]~121_combout ))))

	.dataa(\rfif.rdat2[26]~116_combout ),
	.datab(\rfif.rdat2[26]~123_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[26]~121_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~124_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~124 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[26]~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \rfif.rdat2[26]~106 (
// Equation(s):
// \rfif.rdat2[26]~106_combout  = (\rfif.rdat2[26]~105_combout  & ((\regs[29][26]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[26]~105_combout  & (((\regs[21][26]~q  & Instr_IF_18))))

	.dataa(\rfif.rdat2[26]~105_combout ),
	.datab(\regs[29][26]~q ),
	.datac(\regs[21][26]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~106_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~106 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[26]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[26]~109 (
// Equation(s):
// \rfif.rdat2[26]~109_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][26]~q ))) # (!Instr_IF_18 & (\regs[16][26]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][26]~q ),
	.datad(\regs[20][26]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~109_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~109 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[26]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[26]~110 (
// Equation(s):
// \rfif.rdat2[26]~110_combout  = (Instr_IF_19 & ((\rfif.rdat2[26]~109_combout  & ((\regs[28][26]~q ))) # (!\rfif.rdat2[26]~109_combout  & (\regs[24][26]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[26]~109_combout ))))

	.dataa(\regs[24][26]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[28][26]~q ),
	.datad(\rfif.rdat2[26]~109_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~110_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~110 .lut_mask = 16'hF388;
defparam \rfif.rdat2[26]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \rfif.rdat2[26]~111 (
// Equation(s):
// \rfif.rdat2[26]~111_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\rfif.rdat2[26]~108_combout )) # (!Instr_IF_17 & ((\rfif.rdat2[26]~110_combout )))))

	.dataa(\rfif.rdat2[26]~108_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[26]~110_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~111_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~111 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[26]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[26]~112 (
// Equation(s):
// \rfif.rdat2[26]~112_combout  = (Instr_IF_19 & (((\regs[27][26]~q ) # (Instr_IF_18)))) # (!Instr_IF_19 & (\regs[19][26]~q  & ((!Instr_IF_18))))

	.dataa(\regs[19][26]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[27][26]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~112_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~112 .lut_mask = 16'hCCE2;
defparam \rfif.rdat2[26]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[26]~113 (
// Equation(s):
// \rfif.rdat2[26]~113_combout  = (Instr_IF_18 & ((\rfif.rdat2[26]~112_combout  & ((\regs[31][26]~q ))) # (!\rfif.rdat2[26]~112_combout  & (\regs[23][26]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[26]~112_combout ))))

	.dataa(\regs[23][26]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[31][26]~q ),
	.datad(\rfif.rdat2[26]~112_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~113_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~113 .lut_mask = 16'hF388;
defparam \rfif.rdat2[26]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \rfif.rdat2[26]~114 (
// Equation(s):
// \rfif.rdat2[26]~114_combout  = (Instr_IF_16 & ((\rfif.rdat2[26]~111_combout  & ((\rfif.rdat2[26]~113_combout ))) # (!\rfif.rdat2[26]~111_combout  & (\rfif.rdat2[26]~106_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[26]~111_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[26]~106_combout ),
	.datac(\rfif.rdat2[26]~111_combout ),
	.datad(\rfif.rdat2[26]~113_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[26]~114_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[26]~114 .lut_mask = 16'hF858;
defparam \rfif.rdat2[26]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N25
dffeas \regs[23][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][25] .is_wysiwyg = "true";
defparam \regs[23][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N23
dffeas \regs[19][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][25] .is_wysiwyg = "true";
defparam \regs[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[25]~127 (
// Equation(s):
// \rfif.rdat1[25]~127_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][25]~q )) # (!Instr_IF_23 & ((\regs[19][25]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][25]~q ),
	.datad(\regs[19][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~127_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~127 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[25]~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N11
dffeas \regs[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][25] .is_wysiwyg = "true";
defparam \regs[27][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N1
dffeas \regs[31][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][25] .is_wysiwyg = "true";
defparam \regs[31][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[25]~128 (
// Equation(s):
// \rfif.rdat1[25]~128_combout  = (Instr_IF_24 & ((\rfif.rdat1[25]~127_combout  & ((\regs[31][25]~q ))) # (!\rfif.rdat1[25]~127_combout  & (\regs[27][25]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[25]~127_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[25]~127_combout ),
	.datac(\regs[27][25]~q ),
	.datad(\regs[31][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~128_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~128 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[25]~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N15
dffeas \regs[26][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][25] .is_wysiwyg = "true";
defparam \regs[26][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N19
dffeas \regs[18][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][25] .is_wysiwyg = "true";
defparam \regs[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \rfif.rdat1[25]~120 (
// Equation(s):
// \rfif.rdat1[25]~120_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][25]~q )) # (!Instr_IF_24 & ((\regs[18][25]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][25]~q ),
	.datad(\regs[18][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~120_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~120 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[25]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N13
dffeas \regs[30][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][25] .is_wysiwyg = "true";
defparam \regs[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N25
dffeas \regs[22][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][25] .is_wysiwyg = "true";
defparam \regs[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \rfif.rdat1[25]~121 (
// Equation(s):
// \rfif.rdat1[25]~121_combout  = (Instr_IF_23 & ((\rfif.rdat1[25]~120_combout  & (\regs[30][25]~q )) # (!\rfif.rdat1[25]~120_combout  & ((\regs[22][25]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[25]~120_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[25]~120_combout ),
	.datac(\regs[30][25]~q ),
	.datad(\regs[22][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~121_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~121 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[25]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas \regs[29][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][25] .is_wysiwyg = "true";
defparam \regs[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \regs[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][25] .is_wysiwyg = "true";
defparam \regs[25][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[25]~123 (
// Equation(s):
// \rfif.rdat1[25]~123_combout  = (\rfif.rdat1[25]~122_combout  & ((\regs[29][25]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[25]~122_combout  & (((\regs[25][25]~q  & Instr_IF_24))))

	.dataa(\rfif.rdat1[25]~122_combout ),
	.datab(\regs[29][25]~q ),
	.datac(\regs[25][25]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~123_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~123 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[25]~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N4
cycloneive_lcell_comb \regs[20][25]~feeder (
// Equation(s):
// \regs[20][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b5),
	.cin(gnd),
	.combout(\regs[20][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N5
dffeas \regs[20][25] (
	.clk(!CLK),
	.d(\regs[20][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][25] .is_wysiwyg = "true";
defparam \regs[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N29
dffeas \regs[16][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][25] .is_wysiwyg = "true";
defparam \regs[16][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N27
dffeas \regs[24][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][25] .is_wysiwyg = "true";
defparam \regs[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[25]~124 (
// Equation(s):
// \rfif.rdat1[25]~124_combout  = (Instr_IF_24 & (((\regs[24][25]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[16][25]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[16][25]~q ),
	.datac(\regs[24][25]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~124_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~124 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[25]~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[25]~125 (
// Equation(s):
// \rfif.rdat1[25]~125_combout  = (\rfif.rdat1[25]~124_combout  & ((\regs[28][25]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[25]~124_combout  & (((\regs[20][25]~q  & Instr_IF_23))))

	.dataa(\regs[28][25]~q ),
	.datab(\regs[20][25]~q ),
	.datac(\rfif.rdat1[25]~124_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~125_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~125 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[25]~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[25]~126 (
// Equation(s):
// \rfif.rdat1[25]~126_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\rfif.rdat1[25]~123_combout )) # (!Instr_IF_21 & ((\rfif.rdat1[25]~125_combout )))))

	.dataa(\rfif.rdat1[25]~123_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[25]~125_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~126_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~126 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[25]~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \regs[3][25]~feeder (
// Equation(s):
// \regs[3][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b5),
	.cin(gnd),
	.combout(\regs[3][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N15
dffeas \regs[3][25] (
	.clk(!CLK),
	.d(\regs[3][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][25] .is_wysiwyg = "true";
defparam \regs[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N3
dffeas \regs[2][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][25] .is_wysiwyg = "true";
defparam \regs[2][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N29
dffeas \regs[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][25] .is_wysiwyg = "true";
defparam \regs[1][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N13
dffeas \regs[0][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][25] .is_wysiwyg = "true";
defparam \regs[0][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[25]~134 (
// Equation(s):
// \rfif.rdat1[25]~134_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][25]~q )) # (!Instr_IF_21 & ((\regs[0][25]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][25]~q ),
	.datad(\regs[0][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~134_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~134 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[25]~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[25]~135 (
// Equation(s):
// \rfif.rdat1[25]~135_combout  = (Instr_IF_22 & ((\rfif.rdat1[25]~134_combout  & (\regs[3][25]~q )) # (!\rfif.rdat1[25]~134_combout  & ((\regs[2][25]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[25]~134_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[3][25]~q ),
	.datac(\regs[2][25]~q ),
	.datad(\rfif.rdat1[25]~134_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~135_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~135 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[25]~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \regs[7][25]~feeder (
// Equation(s):
// \regs[7][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b5),
	.cin(gnd),
	.combout(\regs[7][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[7][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N9
dffeas \regs[7][25] (
	.clk(!CLK),
	.d(\regs[7][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][25] .is_wysiwyg = "true";
defparam \regs[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N31
dffeas \regs[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][25] .is_wysiwyg = "true";
defparam \regs[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \rfif.rdat1[25]~133 (
// Equation(s):
// \rfif.rdat1[25]~133_combout  = (\rfif.rdat1[25]~132_combout  & ((\regs[7][25]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[25]~132_combout  & (((\regs[5][25]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[25]~132_combout ),
	.datab(\regs[7][25]~q ),
	.datac(\regs[5][25]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~133_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~133 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[25]~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \rfif.rdat1[25]~136 (
// Equation(s):
// \rfif.rdat1[25]~136_combout  = (Instr_IF_23 & (((Instr_IF_24) # (\rfif.rdat1[25]~133_combout )))) # (!Instr_IF_23 & (\rfif.rdat1[25]~135_combout  & (!Instr_IF_24)))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[25]~135_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[25]~133_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~136_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~136 .lut_mask = 16'hAEA4;
defparam \rfif.rdat1[25]~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N27
dffeas \regs[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][25] .is_wysiwyg = "true";
defparam \regs[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \regs[9][25]~feeder (
// Equation(s):
// \regs[9][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b5),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][25]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N29
dffeas \regs[9][25] (
	.clk(!CLK),
	.d(\regs[9][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][25] .is_wysiwyg = "true";
defparam \regs[9][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \rfif.rdat1[25]~130 (
// Equation(s):
// \rfif.rdat1[25]~130_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][25]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & (\regs[8][25]~q )))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[8][25]~q ),
	.datad(\regs[9][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~130_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~130 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[25]~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N9
dffeas \regs[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][25] .is_wysiwyg = "true";
defparam \regs[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \regs[11][25]~feeder (
// Equation(s):
// \regs[11][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b5),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][25]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N19
dffeas \regs[11][25] (
	.clk(!CLK),
	.d(\regs[11][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][25] .is_wysiwyg = "true";
defparam \regs[11][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[25]~131 (
// Equation(s):
// \rfif.rdat1[25]~131_combout  = (Instr_IF_22 & ((\rfif.rdat1[25]~130_combout  & ((\regs[11][25]~q ))) # (!\rfif.rdat1[25]~130_combout  & (\regs[10][25]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[25]~130_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[25]~130_combout ),
	.datac(\regs[10][25]~q ),
	.datad(\regs[11][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~131_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~131 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[25]~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N16
cycloneive_lcell_comb \regs[15][25]~feeder (
// Equation(s):
// \regs[15][25]~feeder_combout  = \input_b~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b5),
	.cin(gnd),
	.combout(\regs[15][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][25]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N17
dffeas \regs[15][25] (
	.clk(!CLK),
	.d(\regs[15][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][25] .is_wysiwyg = "true";
defparam \regs[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N5
dffeas \regs[12][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][25] .is_wysiwyg = "true";
defparam \regs[12][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N11
dffeas \regs[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][25] .is_wysiwyg = "true";
defparam \regs[14][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \rfif.rdat1[25]~137 (
// Equation(s):
// \rfif.rdat1[25]~137_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[14][25]~q ))) # (!Instr_IF_22 & (\regs[12][25]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][25]~q ),
	.datac(\regs[14][25]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~137_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~137 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[25]~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N21
dffeas \regs[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][25] .is_wysiwyg = "true";
defparam \regs[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \rfif.rdat1[25]~138 (
// Equation(s):
// \rfif.rdat1[25]~138_combout  = (Instr_IF_21 & ((\rfif.rdat1[25]~137_combout  & (\regs[15][25]~q )) # (!\rfif.rdat1[25]~137_combout  & ((\regs[13][25]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[25]~137_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[15][25]~q ),
	.datac(\rfif.rdat1[25]~137_combout ),
	.datad(\regs[13][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[25]~138_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[25]~138 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[25]~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \rfif.rdat2[25]~136 (
// Equation(s):
// \rfif.rdat2[25]~136_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[9][25]~q ))) # (!Instr_IF_16 & (\regs[8][25]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[8][25]~q ),
	.datad(\regs[9][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~136_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~136 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[25]~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \rfif.rdat2[25]~137 (
// Equation(s):
// \rfif.rdat2[25]~137_combout  = (Instr_IF_17 & ((\rfif.rdat2[25]~136_combout  & (\regs[11][25]~q )) # (!\rfif.rdat2[25]~136_combout  & ((\regs[10][25]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[25]~136_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[11][25]~q ),
	.datac(\regs[10][25]~q ),
	.datad(\rfif.rdat2[25]~136_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~137_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~137 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[25]~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \rfif.rdat2[25]~143 (
// Equation(s):
// \rfif.rdat2[25]~143_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][25]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][25]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][25]~q ),
	.datad(\regs[14][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~143_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~143 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[25]~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[25]~144 (
// Equation(s):
// \rfif.rdat2[25]~144_combout  = (Instr_IF_16 & ((\rfif.rdat2[25]~143_combout  & (\regs[15][25]~q )) # (!\rfif.rdat2[25]~143_combout  & ((\regs[13][25]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[25]~143_combout ))))

	.dataa(\regs[15][25]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[13][25]~q ),
	.datad(\rfif.rdat2[25]~143_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~144_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~144 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[25]~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N1
dffeas \regs[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][25] .is_wysiwyg = "true";
defparam \regs[4][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N3
dffeas \regs[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][25] .is_wysiwyg = "true";
defparam \regs[6][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[25]~138 (
// Equation(s):
// \rfif.rdat2[25]~138_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][25]~q ))) # (!Instr_IF_17 & (\regs[4][25]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][25]~q ),
	.datad(\regs[6][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~138_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~138 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[25]~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \rfif.rdat2[25]~139 (
// Equation(s):
// \rfif.rdat2[25]~139_combout  = (Instr_IF_16 & ((\rfif.rdat2[25]~138_combout  & ((\regs[7][25]~q ))) # (!\rfif.rdat2[25]~138_combout  & (\regs[5][25]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[25]~138_combout ))))

	.dataa(\regs[5][25]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[7][25]~q ),
	.datad(\rfif.rdat2[25]~138_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~139_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~139 .lut_mask = 16'hF388;
defparam \rfif.rdat2[25]~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \rfif.rdat2[25]~142 (
// Equation(s):
// \rfif.rdat2[25]~142_combout  = (Instr_IF_18 & (((\rfif.rdat2[25]~139_combout ) # (Instr_IF_19)))) # (!Instr_IF_18 & (\rfif.rdat2[25]~141_combout  & ((!Instr_IF_19))))

	.dataa(\rfif.rdat2[25]~141_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[25]~139_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~142_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~142 .lut_mask = 16'hCCE2;
defparam \rfif.rdat2[25]~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[25]~145 (
// Equation(s):
// \rfif.rdat2[25]~145_combout  = (Instr_IF_19 & ((\rfif.rdat2[25]~142_combout  & ((\rfif.rdat2[25]~144_combout ))) # (!\rfif.rdat2[25]~142_combout  & (\rfif.rdat2[25]~137_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[25]~142_combout ))))

	.dataa(\rfif.rdat2[25]~137_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[25]~144_combout ),
	.datad(\rfif.rdat2[25]~142_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~145_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~145 .lut_mask = 16'hF388;
defparam \rfif.rdat2[25]~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \rfif.rdat2[25]~126 (
// Equation(s):
// \rfif.rdat2[25]~126_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][25]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][25]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][25]~q ),
	.datad(\regs[26][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~126_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~126 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[25]~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[25]~127 (
// Equation(s):
// \rfif.rdat2[25]~127_combout  = (Instr_IF_18 & ((\rfif.rdat2[25]~126_combout  & (\regs[30][25]~q )) # (!\rfif.rdat2[25]~126_combout  & ((\regs[22][25]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[25]~126_combout ))))

	.dataa(\regs[30][25]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][25]~q ),
	.datad(\rfif.rdat2[25]~126_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~127_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~127 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[25]~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[25]~133 (
// Equation(s):
// \rfif.rdat2[25]~133_combout  = (Instr_IF_18 & ((\regs[23][25]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[19][25]~q  & !Instr_IF_19))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][25]~q ),
	.datac(\regs[19][25]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~133_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~133 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[25]~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[25]~134 (
// Equation(s):
// \rfif.rdat2[25]~134_combout  = (\rfif.rdat2[25]~133_combout  & (((\regs[31][25]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[25]~133_combout  & (\regs[27][25]~q  & ((Instr_IF_19))))

	.dataa(\regs[27][25]~q ),
	.datab(\rfif.rdat2[25]~133_combout ),
	.datac(\regs[31][25]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~134_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~134 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[25]~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N23
dffeas \regs[17][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][25] .is_wysiwyg = "true";
defparam \regs[17][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N13
dffeas \regs[21][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][25] .is_wysiwyg = "true";
defparam \regs[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[25]~128 (
// Equation(s):
// \rfif.rdat2[25]~128_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[21][25]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[17][25]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][25]~q ),
	.datad(\regs[21][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~128_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~128 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[25]~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[25]~129 (
// Equation(s):
// \rfif.rdat2[25]~129_combout  = (Instr_IF_19 & ((\rfif.rdat2[25]~128_combout  & ((\regs[29][25]~q ))) # (!\rfif.rdat2[25]~128_combout  & (\regs[25][25]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[25]~128_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][25]~q ),
	.datac(\regs[29][25]~q ),
	.datad(\rfif.rdat2[25]~128_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~129_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~129 .lut_mask = 16'hF588;
defparam \rfif.rdat2[25]~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[25]~130 (
// Equation(s):
// \rfif.rdat2[25]~130_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[24][25]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[16][25]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][25]~q ),
	.datad(\regs[24][25]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~130_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~130 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[25]~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[25]~131 (
// Equation(s):
// \rfif.rdat2[25]~131_combout  = (Instr_IF_18 & ((\rfif.rdat2[25]~130_combout  & (\regs[28][25]~q )) # (!\rfif.rdat2[25]~130_combout  & ((\regs[20][25]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[25]~130_combout ))))

	.dataa(\regs[28][25]~q ),
	.datab(\regs[20][25]~q ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[25]~130_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~131_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~131 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[25]~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \rfif.rdat2[25]~132 (
// Equation(s):
// \rfif.rdat2[25]~132_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[25]~129_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[25]~131_combout )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[25]~129_combout ),
	.datad(\rfif.rdat2[25]~131_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~132_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~132 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[25]~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \rfif.rdat2[25]~135 (
// Equation(s):
// \rfif.rdat2[25]~135_combout  = (Instr_IF_17 & ((\rfif.rdat2[25]~132_combout  & ((\rfif.rdat2[25]~134_combout ))) # (!\rfif.rdat2[25]~132_combout  & (\rfif.rdat2[25]~127_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[25]~132_combout ))))

	.dataa(\rfif.rdat2[25]~127_combout ),
	.datab(\rfif.rdat2[25]~134_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[25]~132_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[25]~135_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[25]~135 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[25]~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N5
dffeas \regs[21][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][24] .is_wysiwyg = "true";
defparam \regs[21][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N7
dffeas \regs[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][24] .is_wysiwyg = "true";
defparam \regs[17][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \regs[25][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][24] .is_wysiwyg = "true";
defparam \regs[25][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[24]~140 (
// Equation(s):
// \rfif.rdat1[24]~140_combout  = (Instr_IF_24 & (((\regs[25][24]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][24]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][24]~q ),
	.datac(\regs[25][24]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~140_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~140 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[24]~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \regs[29][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][24] .is_wysiwyg = "true";
defparam \regs[29][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \rfif.rdat1[24]~141 (
// Equation(s):
// \rfif.rdat1[24]~141_combout  = (\rfif.rdat1[24]~140_combout  & (((\regs[29][24]~q ) # (!Instr_IF_23)))) # (!\rfif.rdat1[24]~140_combout  & (\regs[21][24]~q  & ((Instr_IF_23))))

	.dataa(\regs[21][24]~q ),
	.datab(\rfif.rdat1[24]~140_combout ),
	.datac(\regs[29][24]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~141_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~141 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[24]~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \regs[24][24]~feeder (
// Equation(s):
// \regs[24][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[24][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N5
dffeas \regs[24][24] (
	.clk(!CLK),
	.d(\regs[24][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][24] .is_wysiwyg = "true";
defparam \regs[24][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N27
dffeas \regs[20][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][24] .is_wysiwyg = "true";
defparam \regs[20][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N15
dffeas \regs[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][24] .is_wysiwyg = "true";
defparam \regs[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[24]~144 (
// Equation(s):
// \rfif.rdat1[24]~144_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[20][24]~q )) # (!Instr_IF_23 & ((\regs[16][24]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[20][24]~q ),
	.datad(\regs[16][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~144_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~144 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[24]~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[24]~145 (
// Equation(s):
// \rfif.rdat1[24]~145_combout  = (\rfif.rdat1[24]~144_combout  & ((\regs[28][24]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[24]~144_combout  & (((\regs[24][24]~q  & Instr_IF_24))))

	.dataa(\regs[28][24]~q ),
	.datab(\regs[24][24]~q ),
	.datac(\rfif.rdat1[24]~144_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~145_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~145 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[24]~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N25
dffeas \regs[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][24] .is_wysiwyg = "true";
defparam \regs[26][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N17
dffeas \regs[22][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][24] .is_wysiwyg = "true";
defparam \regs[22][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \rfif.rdat1[24]~142 (
// Equation(s):
// \rfif.rdat1[24]~142_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][24]~q ))) # (!Instr_IF_23 & (\regs[18][24]~q ))))

	.dataa(\regs[18][24]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[22][24]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~142_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~142 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[24]~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[24]~143 (
// Equation(s):
// \rfif.rdat1[24]~143_combout  = (Instr_IF_24 & ((\rfif.rdat1[24]~142_combout  & (\regs[30][24]~q )) # (!\rfif.rdat1[24]~142_combout  & ((\regs[26][24]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[24]~142_combout ))))

	.dataa(\regs[30][24]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[26][24]~q ),
	.datad(\rfif.rdat1[24]~142_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~143_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~143 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[24]~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[24]~146 (
// Equation(s):
// \rfif.rdat1[24]~146_combout  = (Instr_IF_22 & (((Instr_IF_21) # (\rfif.rdat1[24]~143_combout )))) # (!Instr_IF_22 & (\rfif.rdat1[24]~145_combout  & (!Instr_IF_21)))

	.dataa(\rfif.rdat1[24]~145_combout ),
	.datab(Instr_IF_22),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[24]~143_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~146_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~146 .lut_mask = 16'hCEC2;
defparam \rfif.rdat1[24]~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N0
cycloneive_lcell_comb \regs[23][24]~feeder (
// Equation(s):
// \regs[23][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[23][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N1
dffeas \regs[23][24] (
	.clk(!CLK),
	.d(\regs[23][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][24] .is_wysiwyg = "true";
defparam \regs[23][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N30
cycloneive_lcell_comb \regs[27][24]~feeder (
// Equation(s):
// \regs[27][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[27][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N31
dffeas \regs[27][24] (
	.clk(!CLK),
	.d(\regs[27][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][24] .is_wysiwyg = "true";
defparam \regs[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N1
dffeas \regs[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][24] .is_wysiwyg = "true";
defparam \regs[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[24]~147 (
// Equation(s):
// \rfif.rdat1[24]~147_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[27][24]~q )) # (!Instr_IF_24 & ((\regs[19][24]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[27][24]~q ),
	.datad(\regs[19][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~147_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~147 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[24]~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \regs[31][24]~feeder (
// Equation(s):
// \regs[31][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][24]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N1
dffeas \regs[31][24] (
	.clk(!CLK),
	.d(\regs[31][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][24] .is_wysiwyg = "true";
defparam \regs[31][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N22
cycloneive_lcell_comb \rfif.rdat1[24]~148 (
// Equation(s):
// \rfif.rdat1[24]~148_combout  = (Instr_IF_23 & ((\rfif.rdat1[24]~147_combout  & ((\regs[31][24]~q ))) # (!\rfif.rdat1[24]~147_combout  & (\regs[23][24]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[24]~147_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[23][24]~q ),
	.datac(\rfif.rdat1[24]~147_combout ),
	.datad(\regs[31][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~148_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~148 .lut_mask = 16'hF858;
defparam \rfif.rdat1[24]~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \regs[15][24]~feeder (
// Equation(s):
// \regs[15][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[15][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \regs[15][24] (
	.clk(!CLK),
	.d(\regs[15][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][24] .is_wysiwyg = "true";
defparam \regs[15][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \regs[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][24] .is_wysiwyg = "true";
defparam \regs[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \regs[13][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][24] .is_wysiwyg = "true";
defparam \regs[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \rfif.rdat1[24]~157 (
// Equation(s):
// \rfif.rdat1[24]~157_combout  = (Instr_IF_21 & (((\regs[13][24]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][24]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][24]~q ),
	.datac(\regs[13][24]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~157_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~157 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[24]~157 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \regs[14][24]~feeder (
// Equation(s):
// \regs[14][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N11
dffeas \regs[14][24] (
	.clk(!CLK),
	.d(\regs[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][24] .is_wysiwyg = "true";
defparam \regs[14][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \rfif.rdat1[24]~158 (
// Equation(s):
// \rfif.rdat1[24]~158_combout  = (Instr_IF_22 & ((\rfif.rdat1[24]~157_combout  & (\regs[15][24]~q )) # (!\rfif.rdat1[24]~157_combout  & ((\regs[14][24]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[24]~157_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[15][24]~q ),
	.datac(\rfif.rdat1[24]~157_combout ),
	.datad(\regs[14][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~158_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~158 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[24]~158 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N15
dffeas \regs[6][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][24] .is_wysiwyg = "true";
defparam \regs[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N29
dffeas \regs[7][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][24] .is_wysiwyg = "true";
defparam \regs[7][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N7
dffeas \regs[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][24] .is_wysiwyg = "true";
defparam \regs[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[24]~150 (
// Equation(s):
// \rfif.rdat1[24]~150_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][24]~q ))) # (!Instr_IF_21 & (\regs[4][24]~q ))))

	.dataa(\regs[4][24]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][24]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~150_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~150 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[24]~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[24]~151 (
// Equation(s):
// \rfif.rdat1[24]~151_combout  = (Instr_IF_22 & ((\rfif.rdat1[24]~150_combout  & ((\regs[7][24]~q ))) # (!\rfif.rdat1[24]~150_combout  & (\regs[6][24]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[24]~150_combout ))))

	.dataa(\regs[6][24]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[7][24]~q ),
	.datad(\rfif.rdat1[24]~150_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~151_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~151 .lut_mask = 16'hF388;
defparam \rfif.rdat1[24]~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \regs[1][24]~feeder (
// Equation(s):
// \regs[1][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b6),
	.cin(gnd),
	.combout(\regs[1][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][24]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N9
dffeas \regs[1][24] (
	.clk(!CLK),
	.d(\regs[1][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][24] .is_wysiwyg = "true";
defparam \regs[1][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N19
dffeas \regs[2][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][24] .is_wysiwyg = "true";
defparam \regs[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N13
dffeas \regs[0][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][24] .is_wysiwyg = "true";
defparam \regs[0][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[24]~154 (
// Equation(s):
// \rfif.rdat1[24]~154_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][24]~q )) # (!Instr_IF_22 & ((\regs[0][24]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[2][24]~q ),
	.datad(\regs[0][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~154_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~154 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[24]~154 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[24]~155 (
// Equation(s):
// \rfif.rdat1[24]~155_combout  = (Instr_IF_21 & ((\rfif.rdat1[24]~154_combout  & (\regs[3][24]~q )) # (!\rfif.rdat1[24]~154_combout  & ((\regs[1][24]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[24]~154_combout ))))

	.dataa(\regs[3][24]~q ),
	.datab(\regs[1][24]~q ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[24]~154_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~155_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~155 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[24]~155 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N23
dffeas \regs[11][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][24] .is_wysiwyg = "true";
defparam \regs[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N25
dffeas \regs[9][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][24] .is_wysiwyg = "true";
defparam \regs[9][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \regs[10][24]~feeder (
// Equation(s):
// \regs[10][24]~feeder_combout  = \input_b~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][24]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N29
dffeas \regs[10][24] (
	.clk(!CLK),
	.d(\regs[10][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][24] .is_wysiwyg = "true";
defparam \regs[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[24]~152 (
// Equation(s):
// \rfif.rdat1[24]~152_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[10][24]~q ))) # (!Instr_IF_22 & (\regs[8][24]~q ))))

	.dataa(\regs[8][24]~q ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\regs[10][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~152_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~152 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[24]~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[24]~153 (
// Equation(s):
// \rfif.rdat1[24]~153_combout  = (Instr_IF_21 & ((\rfif.rdat1[24]~152_combout  & (\regs[11][24]~q )) # (!\rfif.rdat1[24]~152_combout  & ((\regs[9][24]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[24]~152_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][24]~q ),
	.datac(\regs[9][24]~q ),
	.datad(\rfif.rdat1[24]~152_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~153_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~153 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[24]~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[24]~156 (
// Equation(s):
// \rfif.rdat1[24]~156_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[24]~153_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[24]~155_combout ))))

	.dataa(\rfif.rdat1[24]~155_combout ),
	.datab(Instr_IF_23),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[24]~153_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[24]~156_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[24]~156 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[24]~156 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[24]~147 (
// Equation(s):
// \rfif.rdat2[24]~147_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][24]~q ))) # (!Instr_IF_19 & (\regs[17][24]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][24]~q ),
	.datad(\regs[25][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~147_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~147 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[24]~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \rfif.rdat2[24]~148 (
// Equation(s):
// \rfif.rdat2[24]~148_combout  = (Instr_IF_18 & ((\rfif.rdat2[24]~147_combout  & (\regs[29][24]~q )) # (!\rfif.rdat2[24]~147_combout  & ((\regs[21][24]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[24]~147_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[29][24]~q ),
	.datac(\regs[21][24]~q ),
	.datad(\rfif.rdat2[24]~147_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~148_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~148 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[24]~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \rfif.rdat2[24]~155 (
// Equation(s):
// \rfif.rdat2[24]~155_combout  = (\rfif.rdat2[24]~154_combout  & (((\regs[31][24]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[24]~154_combout  & (\regs[23][24]~q  & (Instr_IF_18)))

	.dataa(\rfif.rdat2[24]~154_combout ),
	.datab(\regs[23][24]~q ),
	.datac(Instr_IF_18),
	.datad(\regs[31][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~155_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~155 .lut_mask = 16'hEA4A;
defparam \rfif.rdat2[24]~155 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N27
dffeas \regs[30][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][24] .is_wysiwyg = "true";
defparam \regs[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N11
dffeas \regs[18][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][24] .is_wysiwyg = "true";
defparam \regs[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \rfif.rdat2[24]~149 (
// Equation(s):
// \rfif.rdat2[24]~149_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][24]~q ))) # (!Instr_IF_18 & (\regs[18][24]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][24]~q ),
	.datad(\regs[22][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~149_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~149 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[24]~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[24]~150 (
// Equation(s):
// \rfif.rdat2[24]~150_combout  = (Instr_IF_19 & ((\rfif.rdat2[24]~149_combout  & ((\regs[30][24]~q ))) # (!\rfif.rdat2[24]~149_combout  & (\regs[26][24]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[24]~149_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][24]~q ),
	.datac(\regs[30][24]~q ),
	.datad(\rfif.rdat2[24]~149_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~150_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~150 .lut_mask = 16'hF588;
defparam \rfif.rdat2[24]~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \rfif.rdat2[24]~153 (
// Equation(s):
// \rfif.rdat2[24]~153_combout  = (Instr_IF_17 & (((Instr_IF_16) # (\rfif.rdat2[24]~150_combout )))) # (!Instr_IF_17 & (\rfif.rdat2[24]~152_combout  & (!Instr_IF_16)))

	.dataa(\rfif.rdat2[24]~152_combout ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[24]~150_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~153_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~153 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[24]~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \rfif.rdat2[24]~156 (
// Equation(s):
// \rfif.rdat2[24]~156_combout  = (Instr_IF_16 & ((\rfif.rdat2[24]~153_combout  & ((\rfif.rdat2[24]~155_combout ))) # (!\rfif.rdat2[24]~153_combout  & (\rfif.rdat2[24]~148_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[24]~153_combout ))))

	.dataa(\rfif.rdat2[24]~148_combout ),
	.datab(\rfif.rdat2[24]~155_combout ),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[24]~153_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~156_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~156 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[24]~156 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \rfif.rdat2[24]~164 (
// Equation(s):
// \rfif.rdat2[24]~164_combout  = (Instr_IF_16 & ((\regs[13][24]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[12][24]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[13][24]~q ),
	.datac(\regs[12][24]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~164_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~164 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[24]~164 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \rfif.rdat2[24]~165 (
// Equation(s):
// \rfif.rdat2[24]~165_combout  = (\rfif.rdat2[24]~164_combout  & (((\regs[15][24]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[24]~164_combout  & (\regs[14][24]~q  & (Instr_IF_17)))

	.dataa(\regs[14][24]~q ),
	.datab(\rfif.rdat2[24]~164_combout ),
	.datac(Instr_IF_17),
	.datad(\regs[15][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~165_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~165 .lut_mask = 16'hEC2C;
defparam \rfif.rdat2[24]~165 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[24]~161 (
// Equation(s):
// \rfif.rdat2[24]~161_combout  = (Instr_IF_17 & ((\regs[2][24]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((!Instr_IF_16 & \regs[0][24]~q ))))

	.dataa(Instr_IF_17),
	.datab(\regs[2][24]~q ),
	.datac(Instr_IF_16),
	.datad(\regs[0][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~161_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~161 .lut_mask = 16'hADA8;
defparam \rfif.rdat2[24]~161 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[24]~162 (
// Equation(s):
// \rfif.rdat2[24]~162_combout  = (Instr_IF_16 & ((\rfif.rdat2[24]~161_combout  & (\regs[3][24]~q )) # (!\rfif.rdat2[24]~161_combout  & ((\regs[1][24]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[24]~161_combout ))))

	.dataa(\regs[3][24]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[1][24]~q ),
	.datad(\rfif.rdat2[24]~161_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~162_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~162 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[24]~162 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \rfif.rdat2[24]~163 (
// Equation(s):
// \rfif.rdat2[24]~163_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[24]~160_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[24]~162_combout )))))

	.dataa(\rfif.rdat2[24]~160_combout ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[24]~162_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~163_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~163 .lut_mask = 16'hE3E0;
defparam \rfif.rdat2[24]~163 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N29
dffeas \regs[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][24] .is_wysiwyg = "true";
defparam \regs[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[24]~157 (
// Equation(s):
// \rfif.rdat2[24]~157_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][24]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][24]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][24]~q ),
	.datad(\regs[5][24]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~157_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~157 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[24]~157 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \rfif.rdat2[24]~158 (
// Equation(s):
// \rfif.rdat2[24]~158_combout  = (Instr_IF_17 & ((\rfif.rdat2[24]~157_combout  & (\regs[7][24]~q )) # (!\rfif.rdat2[24]~157_combout  & ((\regs[6][24]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[24]~157_combout ))))

	.dataa(\regs[7][24]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[6][24]~q ),
	.datad(\rfif.rdat2[24]~157_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~158_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~158 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[24]~158 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \rfif.rdat2[24]~166 (
// Equation(s):
// \rfif.rdat2[24]~166_combout  = (Instr_IF_18 & ((\rfif.rdat2[24]~163_combout  & (\rfif.rdat2[24]~165_combout )) # (!\rfif.rdat2[24]~163_combout  & ((\rfif.rdat2[24]~158_combout ))))) # (!Instr_IF_18 & (((\rfif.rdat2[24]~163_combout ))))

	.dataa(\rfif.rdat2[24]~165_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[24]~163_combout ),
	.datad(\rfif.rdat2[24]~158_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[24]~166_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[24]~166 .lut_mask = 16'hBCB0;
defparam \rfif.rdat2[24]~166 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N23
dffeas \regs[26][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][23] .is_wysiwyg = "true";
defparam \regs[26][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N27
dffeas \regs[18][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][23] .is_wysiwyg = "true";
defparam \regs[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \rfif.rdat1[23]~160 (
// Equation(s):
// \rfif.rdat1[23]~160_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][23]~q )) # (!Instr_IF_24 & ((\regs[18][23]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][23]~q ),
	.datad(\regs[18][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~160_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~160 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[23]~160 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N25
dffeas \regs[22][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][23] .is_wysiwyg = "true";
defparam \regs[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N9
dffeas \regs[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][23] .is_wysiwyg = "true";
defparam \regs[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[23]~161 (
// Equation(s):
// \rfif.rdat1[23]~161_combout  = (\rfif.rdat1[23]~160_combout  & (((\regs[30][23]~q ) # (!Instr_IF_23)))) # (!\rfif.rdat1[23]~160_combout  & (\regs[22][23]~q  & ((Instr_IF_23))))

	.dataa(\rfif.rdat1[23]~160_combout ),
	.datab(\regs[22][23]~q ),
	.datac(\regs[30][23]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~161_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~161 .lut_mask = 16'hE4AA;
defparam \rfif.rdat1[23]~161 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N3
dffeas \regs[19][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][23] .is_wysiwyg = "true";
defparam \regs[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N18
cycloneive_lcell_comb \regs[23][23]~feeder (
// Equation(s):
// \regs[23][23]~feeder_combout  = \input_b~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b7),
	.cin(gnd),
	.combout(\regs[23][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][23]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N19
dffeas \regs[23][23] (
	.clk(!CLK),
	.d(\regs[23][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][23] .is_wysiwyg = "true";
defparam \regs[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[23]~167 (
// Equation(s):
// \rfif.rdat1[23]~167_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[23][23]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[19][23]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[19][23]~q ),
	.datad(\regs[23][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~167_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~167 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[23]~167 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N29
dffeas \regs[31][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][23] .is_wysiwyg = "true";
defparam \regs[31][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N31
dffeas \regs[27][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][23] .is_wysiwyg = "true";
defparam \regs[27][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N30
cycloneive_lcell_comb \rfif.rdat1[23]~168 (
// Equation(s):
// \rfif.rdat1[23]~168_combout  = (\rfif.rdat1[23]~167_combout  & ((\regs[31][23]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[23]~167_combout  & (((\regs[27][23]~q  & Instr_IF_24))))

	.dataa(\rfif.rdat1[23]~167_combout ),
	.datab(\regs[31][23]~q ),
	.datac(\regs[27][23]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~168_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~168 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[23]~168 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \regs[25][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][23] .is_wysiwyg = "true";
defparam \regs[25][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N1
dffeas \regs[21][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][23] .is_wysiwyg = "true";
defparam \regs[21][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N3
dffeas \regs[17][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][23] .is_wysiwyg = "true";
defparam \regs[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[23]~162 (
// Equation(s):
// \rfif.rdat1[23]~162_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][23]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & ((\regs[17][23]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[21][23]~q ),
	.datad(\regs[17][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~162_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~162 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[23]~162 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[23]~163 (
// Equation(s):
// \rfif.rdat1[23]~163_combout  = (Instr_IF_24 & ((\rfif.rdat1[23]~162_combout  & (\regs[29][23]~q )) # (!\rfif.rdat1[23]~162_combout  & ((\regs[25][23]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[23]~162_combout ))))

	.dataa(\regs[29][23]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[25][23]~q ),
	.datad(\rfif.rdat1[23]~162_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~163_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~163 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[23]~163 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N21
dffeas \regs[20][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][23] .is_wysiwyg = "true";
defparam \regs[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \regs[24][23]~feeder (
// Equation(s):
// \regs[24][23]~feeder_combout  = \input_b~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][23]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N13
dffeas \regs[24][23] (
	.clk(!CLK),
	.d(\regs[24][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][23] .is_wysiwyg = "true";
defparam \regs[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N19
dffeas \regs[16][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][23] .is_wysiwyg = "true";
defparam \regs[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[23]~164 (
// Equation(s):
// \rfif.rdat1[23]~164_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[24][23]~q )) # (!Instr_IF_24 & ((\regs[16][23]~q )))))

	.dataa(Instr_IF_23),
	.datab(\regs[24][23]~q ),
	.datac(\regs[16][23]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~164_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~164 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[23]~164 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[23]~165 (
// Equation(s):
// \rfif.rdat1[23]~165_combout  = (Instr_IF_23 & ((\rfif.rdat1[23]~164_combout  & (\regs[28][23]~q )) # (!\rfif.rdat1[23]~164_combout  & ((\regs[20][23]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[23]~164_combout ))))

	.dataa(\regs[28][23]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][23]~q ),
	.datad(\rfif.rdat1[23]~164_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~165_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~165 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[23]~165 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[23]~166 (
// Equation(s):
// \rfif.rdat1[23]~166_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\rfif.rdat1[23]~163_combout )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\rfif.rdat1[23]~165_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[23]~163_combout ),
	.datad(\rfif.rdat1[23]~165_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~166_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~166 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[23]~166 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N11
dffeas \regs[0][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][23] .is_wysiwyg = "true";
defparam \regs[0][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \regs[1][23]~feeder (
// Equation(s):
// \regs[1][23]~feeder_combout  = \input_b~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[1][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][23]~feeder .lut_mask = 16'hF0F0;
defparam \regs[1][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N13
dffeas \regs[1][23] (
	.clk(!CLK),
	.d(\regs[1][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][23] .is_wysiwyg = "true";
defparam \regs[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[23]~174 (
// Equation(s):
// \rfif.rdat1[23]~174_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[1][23]~q ))) # (!Instr_IF_21 & (\regs[0][23]~q ))))

	.dataa(Instr_IF_22),
	.datab(\regs[0][23]~q ),
	.datac(Instr_IF_21),
	.datad(\regs[1][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~174_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~174 .lut_mask = 16'hF4A4;
defparam \rfif.rdat1[23]~174 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N25
dffeas \regs[3][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][23] .is_wysiwyg = "true";
defparam \regs[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N9
dffeas \regs[2][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][23] .is_wysiwyg = "true";
defparam \regs[2][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[23]~175 (
// Equation(s):
// \rfif.rdat1[23]~175_combout  = (Instr_IF_22 & ((\rfif.rdat1[23]~174_combout  & (\regs[3][23]~q )) # (!\rfif.rdat1[23]~174_combout  & ((\regs[2][23]~q ))))) # (!Instr_IF_22 & (\rfif.rdat1[23]~174_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[23]~174_combout ),
	.datac(\regs[3][23]~q ),
	.datad(\regs[2][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~175_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~175 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[23]~175 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N17
dffeas \regs[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][23] .is_wysiwyg = "true";
defparam \regs[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N1
dffeas \regs[6][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][23] .is_wysiwyg = "true";
defparam \regs[6][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[23]~172 (
// Equation(s):
// \rfif.rdat1[23]~172_combout  = (Instr_IF_22 & (((\regs[6][23]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[4][23]~q  & ((!Instr_IF_21))))

	.dataa(\regs[4][23]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[6][23]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~172_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~172 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[23]~172 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \rfif.rdat1[23]~173 (
// Equation(s):
// \rfif.rdat1[23]~173_combout  = (Instr_IF_21 & ((\rfif.rdat1[23]~172_combout  & (\regs[7][23]~q )) # (!\rfif.rdat1[23]~172_combout  & ((\regs[5][23]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[23]~172_combout ))))

	.dataa(\regs[7][23]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][23]~q ),
	.datad(\rfif.rdat1[23]~172_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~173_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~173 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[23]~173 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \rfif.rdat1[23]~176 (
// Equation(s):
// \rfif.rdat1[23]~176_combout  = (Instr_IF_23 & (((Instr_IF_24) # (\rfif.rdat1[23]~173_combout )))) # (!Instr_IF_23 & (\rfif.rdat1[23]~175_combout  & (!Instr_IF_24)))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[23]~175_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[23]~173_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~176_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~176 .lut_mask = 16'hAEA4;
defparam \rfif.rdat1[23]~176 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N3
dffeas \regs[14][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][23] .is_wysiwyg = "true";
defparam \regs[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N25
dffeas \regs[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][23] .is_wysiwyg = "true";
defparam \regs[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \rfif.rdat1[23]~177 (
// Equation(s):
// \rfif.rdat1[23]~177_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][23]~q )) # (!Instr_IF_22 & ((\regs[12][23]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[14][23]~q ),
	.datad(\regs[12][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~177_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~177 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[23]~177 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N9
dffeas \regs[15][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][23] .is_wysiwyg = "true";
defparam \regs[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N29
dffeas \regs[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][23] .is_wysiwyg = "true";
defparam \regs[13][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[23]~178 (
// Equation(s):
// \rfif.rdat1[23]~178_combout  = (Instr_IF_21 & ((\rfif.rdat1[23]~177_combout  & (\regs[15][23]~q )) # (!\rfif.rdat1[23]~177_combout  & ((\regs[13][23]~q ))))) # (!Instr_IF_21 & (\rfif.rdat1[23]~177_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[23]~177_combout ),
	.datac(\regs[15][23]~q ),
	.datad(\regs[13][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~178_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~178 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[23]~178 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N15
dffeas \regs[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][23] .is_wysiwyg = "true";
defparam \regs[10][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N17
dffeas \regs[9][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][23] .is_wysiwyg = "true";
defparam \regs[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N13
dffeas \regs[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][23] .is_wysiwyg = "true";
defparam \regs[8][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \rfif.rdat1[23]~170 (
// Equation(s):
// \rfif.rdat1[23]~170_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][23]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[8][23]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[9][23]~q ),
	.datad(\regs[8][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~170_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~170 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[23]~170 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N7
dffeas \regs[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][23] .is_wysiwyg = "true";
defparam \regs[11][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \rfif.rdat1[23]~171 (
// Equation(s):
// \rfif.rdat1[23]~171_combout  = (\rfif.rdat1[23]~170_combout  & (((\regs[11][23]~q ) # (!Instr_IF_22)))) # (!\rfif.rdat1[23]~170_combout  & (\regs[10][23]~q  & ((Instr_IF_22))))

	.dataa(\regs[10][23]~q ),
	.datab(\rfif.rdat1[23]~170_combout ),
	.datac(\regs[11][23]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[23]~171_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[23]~171 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[23]~171 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \rfif.rdat2[23]~179 (
// Equation(s):
// \rfif.rdat2[23]~179_combout  = (\rfif.rdat2[23]~178_combout  & (((\regs[11][23]~q )) # (!Instr_IF_17))) # (!\rfif.rdat2[23]~178_combout  & (Instr_IF_17 & (\regs[10][23]~q )))

	.dataa(\rfif.rdat2[23]~178_combout ),
	.datab(Instr_IF_17),
	.datac(\regs[10][23]~q ),
	.datad(\regs[11][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~179_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~179 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[23]~179 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[23]~185 (
// Equation(s):
// \rfif.rdat2[23]~185_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][23]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][23]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][23]~q ),
	.datad(\regs[14][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~185_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~185 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[23]~185 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \rfif.rdat2[23]~186 (
// Equation(s):
// \rfif.rdat2[23]~186_combout  = (Instr_IF_16 & ((\rfif.rdat2[23]~185_combout  & ((\regs[15][23]~q ))) # (!\rfif.rdat2[23]~185_combout  & (\regs[13][23]~q )))) # (!Instr_IF_16 & (\rfif.rdat2[23]~185_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[23]~185_combout ),
	.datac(\regs[13][23]~q ),
	.datad(\regs[15][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~186_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~186 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[23]~186 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[23]~182 (
// Equation(s):
// \rfif.rdat2[23]~182_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[1][23]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[0][23]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][23]~q ),
	.datad(\regs[1][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~182_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~182 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[23]~182 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[23]~183 (
// Equation(s):
// \rfif.rdat2[23]~183_combout  = (Instr_IF_17 & ((\rfif.rdat2[23]~182_combout  & (\regs[3][23]~q )) # (!\rfif.rdat2[23]~182_combout  & ((\regs[2][23]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[23]~182_combout ))))

	.dataa(\regs[3][23]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[2][23]~q ),
	.datad(\rfif.rdat2[23]~182_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~183_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~183 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[23]~183 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N27
dffeas \regs[7][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][23] .is_wysiwyg = "true";
defparam \regs[7][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[23]~181 (
// Equation(s):
// \rfif.rdat2[23]~181_combout  = (\rfif.rdat2[23]~180_combout  & (((\regs[7][23]~q )) # (!Instr_IF_16))) # (!\rfif.rdat2[23]~180_combout  & (Instr_IF_16 & ((\regs[5][23]~q ))))

	.dataa(\rfif.rdat2[23]~180_combout ),
	.datab(Instr_IF_16),
	.datac(\regs[7][23]~q ),
	.datad(\regs[5][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~181_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~181 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[23]~181 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[23]~184 (
// Equation(s):
// \rfif.rdat2[23]~184_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & ((\rfif.rdat2[23]~181_combout ))) # (!Instr_IF_18 & (\rfif.rdat2[23]~183_combout ))))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[23]~183_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[23]~181_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~184_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~184 .lut_mask = 16'hF4A4;
defparam \rfif.rdat2[23]~184 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \rfif.rdat2[23]~187 (
// Equation(s):
// \rfif.rdat2[23]~187_combout  = (Instr_IF_19 & ((\rfif.rdat2[23]~184_combout  & ((\rfif.rdat2[23]~186_combout ))) # (!\rfif.rdat2[23]~184_combout  & (\rfif.rdat2[23]~179_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[23]~184_combout ))))

	.dataa(\rfif.rdat2[23]~179_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[23]~186_combout ),
	.datad(\rfif.rdat2[23]~184_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~187_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~187 .lut_mask = 16'hF388;
defparam \rfif.rdat2[23]~187 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[23]~169 (
// Equation(s):
// \rfif.rdat2[23]~169_combout  = (\rfif.rdat2[23]~168_combout  & ((\regs[30][23]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[23]~168_combout  & (((\regs[22][23]~q  & Instr_IF_18))))

	.dataa(\rfif.rdat2[23]~168_combout ),
	.datab(\regs[30][23]~q ),
	.datac(\regs[22][23]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~169_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~169 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[23]~169 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[23]~175 (
// Equation(s):
// \rfif.rdat2[23]~175_combout  = (Instr_IF_18 & ((\regs[23][23]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[19][23]~q  & !Instr_IF_19))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][23]~q ),
	.datac(\regs[19][23]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~175_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~175 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[23]~175 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[23]~176 (
// Equation(s):
// \rfif.rdat2[23]~176_combout  = (Instr_IF_19 & ((\rfif.rdat2[23]~175_combout  & ((\regs[31][23]~q ))) # (!\rfif.rdat2[23]~175_combout  & (\regs[27][23]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[23]~175_combout ))))

	.dataa(\regs[27][23]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[31][23]~q ),
	.datad(\rfif.rdat2[23]~175_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~176_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~176 .lut_mask = 16'hF388;
defparam \rfif.rdat2[23]~176 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \regs[29][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][23] .is_wysiwyg = "true";
defparam \regs[29][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \rfif.rdat2[23]~170 (
// Equation(s):
// \rfif.rdat2[23]~170_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[21][23]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[17][23]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][23]~q ),
	.datad(\regs[21][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~170_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~170 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[23]~170 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[23]~171 (
// Equation(s):
// \rfif.rdat2[23]~171_combout  = (Instr_IF_19 & ((\rfif.rdat2[23]~170_combout  & ((\regs[29][23]~q ))) # (!\rfif.rdat2[23]~170_combout  & (\regs[25][23]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[23]~170_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][23]~q ),
	.datac(\regs[29][23]~q ),
	.datad(\rfif.rdat2[23]~170_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~171_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~171 .lut_mask = 16'hF588;
defparam \rfif.rdat2[23]~171 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[23]~172 (
// Equation(s):
// \rfif.rdat2[23]~172_combout  = (Instr_IF_19 & (((Instr_IF_18) # (\regs[24][23]~q )))) # (!Instr_IF_19 & (\regs[16][23]~q  & (!Instr_IF_18)))

	.dataa(Instr_IF_19),
	.datab(\regs[16][23]~q ),
	.datac(Instr_IF_18),
	.datad(\regs[24][23]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~172_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~172 .lut_mask = 16'hAEA4;
defparam \rfif.rdat2[23]~172 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[23]~173 (
// Equation(s):
// \rfif.rdat2[23]~173_combout  = (Instr_IF_18 & ((\rfif.rdat2[23]~172_combout  & (\regs[28][23]~q )) # (!\rfif.rdat2[23]~172_combout  & ((\regs[20][23]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[23]~172_combout ))))

	.dataa(\regs[28][23]~q ),
	.datab(\regs[20][23]~q ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[23]~172_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~173_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~173 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[23]~173 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \rfif.rdat2[23]~174 (
// Equation(s):
// \rfif.rdat2[23]~174_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[23]~171_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[23]~173_combout )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[23]~171_combout ),
	.datad(\rfif.rdat2[23]~173_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~174_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~174 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[23]~174 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[23]~177 (
// Equation(s):
// \rfif.rdat2[23]~177_combout  = (Instr_IF_17 & ((\rfif.rdat2[23]~174_combout  & ((\rfif.rdat2[23]~176_combout ))) # (!\rfif.rdat2[23]~174_combout  & (\rfif.rdat2[23]~169_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[23]~174_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[23]~169_combout ),
	.datac(\rfif.rdat2[23]~176_combout ),
	.datad(\rfif.rdat2[23]~174_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[23]~177_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[23]~177 .lut_mask = 16'hF588;
defparam \rfif.rdat2[23]~177 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \regs[24][22]~feeder (
// Equation(s):
// \regs[24][22]~feeder_combout  = \input_b~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b8),
	.cin(gnd),
	.combout(\regs[24][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[24][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N3
dffeas \regs[24][22] (
	.clk(!CLK),
	.d(\regs[24][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][22] .is_wysiwyg = "true";
defparam \regs[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \regs[28][22]~feeder (
// Equation(s):
// \regs[28][22]~feeder_combout  = \input_b~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b8),
	.cin(gnd),
	.combout(\regs[28][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][22]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N25
dffeas \regs[28][22] (
	.clk(!CLK),
	.d(\regs[28][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][22] .is_wysiwyg = "true";
defparam \regs[28][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[22]~185 (
// Equation(s):
// \rfif.rdat1[22]~185_combout  = (\rfif.rdat1[22]~184_combout  & (((\regs[28][22]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[22]~184_combout  & (Instr_IF_24 & (\regs[24][22]~q )))

	.dataa(\rfif.rdat1[22]~184_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[24][22]~q ),
	.datad(\regs[28][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~185_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~185 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[22]~185 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N1
dffeas \regs[22][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][22] .is_wysiwyg = "true";
defparam \regs[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N11
dffeas \regs[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][22] .is_wysiwyg = "true";
defparam \regs[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[22]~182 (
// Equation(s):
// \rfif.rdat1[22]~182_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[22][22]~q )) # (!Instr_IF_23 & ((\regs[18][22]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[22][22]~q ),
	.datad(\regs[18][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~182_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~182 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[22]~182 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N25
dffeas \regs[26][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][22] .is_wysiwyg = "true";
defparam \regs[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \rfif.rdat1[22]~183 (
// Equation(s):
// \rfif.rdat1[22]~183_combout  = (\rfif.rdat1[22]~182_combout  & ((\regs[30][22]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[22]~182_combout  & (((\regs[26][22]~q  & Instr_IF_24))))

	.dataa(\regs[30][22]~q ),
	.datab(\rfif.rdat1[22]~182_combout ),
	.datac(\regs[26][22]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~183_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~183 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[22]~183 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[22]~186 (
// Equation(s):
// \rfif.rdat1[22]~186_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[22]~183_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[22]~185_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[22]~185_combout ),
	.datad(\rfif.rdat1[22]~183_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~186_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~186 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[22]~186 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N15
dffeas \regs[17][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][22] .is_wysiwyg = "true";
defparam \regs[17][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \regs[25][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][22] .is_wysiwyg = "true";
defparam \regs[25][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[22]~180 (
// Equation(s):
// \rfif.rdat1[22]~180_combout  = (Instr_IF_24 & (((\regs[25][22]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][22]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][22]~q ),
	.datac(\regs[25][22]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~180_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~180 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[22]~180 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \regs[29][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][22] .is_wysiwyg = "true";
defparam \regs[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N5
dffeas \regs[21][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][22] .is_wysiwyg = "true";
defparam \regs[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[22]~181 (
// Equation(s):
// \rfif.rdat1[22]~181_combout  = (Instr_IF_23 & ((\rfif.rdat1[22]~180_combout  & (\regs[29][22]~q )) # (!\rfif.rdat1[22]~180_combout  & ((\regs[21][22]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[22]~180_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[22]~180_combout ),
	.datac(\regs[29][22]~q ),
	.datad(\regs[21][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~181_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~181 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[22]~181 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N12
cycloneive_lcell_comb \regs[23][22]~feeder (
// Equation(s):
// \regs[23][22]~feeder_combout  = \input_b~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N13
dffeas \regs[23][22] (
	.clk(!CLK),
	.d(\regs[23][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][22] .is_wysiwyg = "true";
defparam \regs[23][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N15
dffeas \regs[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][22] .is_wysiwyg = "true";
defparam \regs[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N3
dffeas \regs[27][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][22] .is_wysiwyg = "true";
defparam \regs[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N29
dffeas \regs[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][22] .is_wysiwyg = "true";
defparam \regs[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[22]~187 (
// Equation(s):
// \rfif.rdat1[22]~187_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][22]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][22]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][22]~q ),
	.datad(\regs[19][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~187_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~187 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[22]~187 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N2
cycloneive_lcell_comb \rfif.rdat1[22]~188 (
// Equation(s):
// \rfif.rdat1[22]~188_combout  = (Instr_IF_23 & ((\rfif.rdat1[22]~187_combout  & ((\regs[31][22]~q ))) # (!\rfif.rdat1[22]~187_combout  & (\regs[23][22]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[22]~187_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[23][22]~q ),
	.datac(\regs[31][22]~q ),
	.datad(\rfif.rdat1[22]~187_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~188_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~188 .lut_mask = 16'hF588;
defparam \rfif.rdat1[22]~188 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \regs[14][22]~feeder (
// Equation(s):
// \regs[14][22]~feeder_combout  = \input_b~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N15
dffeas \regs[14][22] (
	.clk(!CLK),
	.d(\regs[14][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][22] .is_wysiwyg = "true";
defparam \regs[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N21
dffeas \regs[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][22] .is_wysiwyg = "true";
defparam \regs[12][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N17
dffeas \regs[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][22] .is_wysiwyg = "true";
defparam \regs[13][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \rfif.rdat1[22]~197 (
// Equation(s):
// \rfif.rdat1[22]~197_combout  = (Instr_IF_21 & (((\regs[13][22]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][22]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][22]~q ),
	.datac(\regs[13][22]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~197_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~197 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[22]~197 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N3
dffeas \regs[15][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][22] .is_wysiwyg = "true";
defparam \regs[15][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \rfif.rdat1[22]~198 (
// Equation(s):
// \rfif.rdat1[22]~198_combout  = (Instr_IF_22 & ((\rfif.rdat1[22]~197_combout  & ((\regs[15][22]~q ))) # (!\rfif.rdat1[22]~197_combout  & (\regs[14][22]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[22]~197_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[14][22]~q ),
	.datac(\rfif.rdat1[22]~197_combout ),
	.datad(\regs[15][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~198_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~198 .lut_mask = 16'hF858;
defparam \rfif.rdat1[22]~198 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \regs[3][22]~feeder (
// Equation(s):
// \regs[3][22]~feeder_combout  = \input_b~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][22]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N17
dffeas \regs[3][22] (
	.clk(!CLK),
	.d(\regs[3][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][22] .is_wysiwyg = "true";
defparam \regs[3][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N3
dffeas \regs[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][22] .is_wysiwyg = "true";
defparam \regs[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N21
dffeas \regs[0][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][22] .is_wysiwyg = "true";
defparam \regs[0][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[22]~194 (
// Equation(s):
// \rfif.rdat1[22]~194_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][22]~q )) # (!Instr_IF_22 & ((\regs[0][22]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[2][22]~q ),
	.datad(\regs[0][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~194_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~194 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[22]~194 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[22]~195 (
// Equation(s):
// \rfif.rdat1[22]~195_combout  = (\rfif.rdat1[22]~194_combout  & (((\regs[3][22]~q ) # (!Instr_IF_21)))) # (!\rfif.rdat1[22]~194_combout  & (\regs[1][22]~q  & ((Instr_IF_21))))

	.dataa(\regs[1][22]~q ),
	.datab(\regs[3][22]~q ),
	.datac(\rfif.rdat1[22]~194_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~195_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~195 .lut_mask = 16'hCAF0;
defparam \rfif.rdat1[22]~195 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N7
dffeas \regs[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][22] .is_wysiwyg = "true";
defparam \regs[10][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N17
dffeas \regs[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][22] .is_wysiwyg = "true";
defparam \regs[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N6
cycloneive_lcell_comb \rfif.rdat1[22]~192 (
// Equation(s):
// \rfif.rdat1[22]~192_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][22]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][22]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][22]~q ),
	.datad(\regs[8][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~192_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~192 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[22]~192 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N21
dffeas \regs[9][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][22] .is_wysiwyg = "true";
defparam \regs[9][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[22]~193 (
// Equation(s):
// \rfif.rdat1[22]~193_combout  = (\rfif.rdat1[22]~192_combout  & ((\regs[11][22]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[22]~192_combout  & (((\regs[9][22]~q  & Instr_IF_21))))

	.dataa(\regs[11][22]~q ),
	.datab(\rfif.rdat1[22]~192_combout ),
	.datac(\regs[9][22]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~193_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~193 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[22]~193 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[22]~196 (
// Equation(s):
// \rfif.rdat1[22]~196_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[22]~193_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[22]~195_combout ))))

	.dataa(\rfif.rdat1[22]~195_combout ),
	.datab(Instr_IF_23),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[22]~193_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~196_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~196 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[22]~196 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N25
dffeas \regs[6][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][22] .is_wysiwyg = "true";
defparam \regs[6][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N9
dffeas \regs[7][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][22] .is_wysiwyg = "true";
defparam \regs[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \regs[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][22] .is_wysiwyg = "true";
defparam \regs[5][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N23
dffeas \regs[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][22] .is_wysiwyg = "true";
defparam \regs[4][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \rfif.rdat1[22]~190 (
// Equation(s):
// \rfif.rdat1[22]~190_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[5][22]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[4][22]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[5][22]~q ),
	.datad(\regs[4][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~190_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~190 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[22]~190 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[22]~191 (
// Equation(s):
// \rfif.rdat1[22]~191_combout  = (Instr_IF_22 & ((\rfif.rdat1[22]~190_combout  & ((\regs[7][22]~q ))) # (!\rfif.rdat1[22]~190_combout  & (\regs[6][22]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[22]~190_combout ))))

	.dataa(\regs[6][22]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[7][22]~q ),
	.datad(\rfif.rdat1[22]~190_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[22]~191_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[22]~191 .lut_mask = 16'hF388;
defparam \rfif.rdat1[22]~191 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N14
cycloneive_lcell_comb \rfif.rdat2[22]~189 (
// Equation(s):
// \rfif.rdat2[22]~189_combout  = (Instr_IF_19 & ((\regs[25][22]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[17][22]~q  & !Instr_IF_18))))

	.dataa(\regs[25][22]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[17][22]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~189_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~189 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[22]~189 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N4
cycloneive_lcell_comb \rfif.rdat2[22]~190 (
// Equation(s):
// \rfif.rdat2[22]~190_combout  = (\rfif.rdat2[22]~189_combout  & ((\regs[29][22]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[22]~189_combout  & (((\regs[21][22]~q  & Instr_IF_18))))

	.dataa(\regs[29][22]~q ),
	.datab(\rfif.rdat2[22]~189_combout ),
	.datac(\regs[21][22]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~190_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~190 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[22]~190 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[22]~196 (
// Equation(s):
// \rfif.rdat2[22]~196_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\regs[27][22]~q )) # (!Instr_IF_19 & ((\regs[19][22]~q )))))

	.dataa(\regs[27][22]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[19][22]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~196_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~196 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[22]~196 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N14
cycloneive_lcell_comb \rfif.rdat2[22]~197 (
// Equation(s):
// \rfif.rdat2[22]~197_combout  = (\rfif.rdat2[22]~196_combout  & (((\regs[31][22]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[22]~196_combout  & (\regs[23][22]~q  & ((Instr_IF_18))))

	.dataa(\regs[23][22]~q ),
	.datab(\rfif.rdat2[22]~196_combout ),
	.datac(\regs[31][22]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~197_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~197 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[22]~197 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N11
dffeas \regs[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][22] .is_wysiwyg = "true";
defparam \regs[16][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \regs[20][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][22] .is_wysiwyg = "true";
defparam \regs[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[22]~193 (
// Equation(s):
// \rfif.rdat2[22]~193_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][22]~q ))) # (!Instr_IF_18 & (\regs[16][22]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][22]~q ),
	.datad(\regs[20][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~193_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~193 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[22]~193 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[22]~194 (
// Equation(s):
// \rfif.rdat2[22]~194_combout  = (Instr_IF_19 & ((\rfif.rdat2[22]~193_combout  & (\regs[28][22]~q )) # (!\rfif.rdat2[22]~193_combout  & ((\regs[24][22]~q ))))) # (!Instr_IF_19 & (((\rfif.rdat2[22]~193_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[28][22]~q ),
	.datac(\rfif.rdat2[22]~193_combout ),
	.datad(\regs[24][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~194_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~194 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[22]~194 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N23
dffeas \regs[30][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][22] .is_wysiwyg = "true";
defparam \regs[30][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \rfif.rdat2[22]~191 (
// Equation(s):
// \rfif.rdat2[22]~191_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][22]~q ))) # (!Instr_IF_18 & (\regs[18][22]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][22]~q ),
	.datad(\regs[22][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~191_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~191 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[22]~191 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \rfif.rdat2[22]~192 (
// Equation(s):
// \rfif.rdat2[22]~192_combout  = (Instr_IF_19 & ((\rfif.rdat2[22]~191_combout  & ((\regs[30][22]~q ))) # (!\rfif.rdat2[22]~191_combout  & (\regs[26][22]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[22]~191_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][22]~q ),
	.datac(\regs[30][22]~q ),
	.datad(\rfif.rdat2[22]~191_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~192_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~192 .lut_mask = 16'hF588;
defparam \rfif.rdat2[22]~192 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[22]~195 (
// Equation(s):
// \rfif.rdat2[22]~195_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[22]~192_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[22]~194_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[22]~194_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[22]~192_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~195_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~195 .lut_mask = 16'hF4A4;
defparam \rfif.rdat2[22]~195 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \rfif.rdat2[22]~198 (
// Equation(s):
// \rfif.rdat2[22]~198_combout  = (Instr_IF_16 & ((\rfif.rdat2[22]~195_combout  & ((\rfif.rdat2[22]~197_combout ))) # (!\rfif.rdat2[22]~195_combout  & (\rfif.rdat2[22]~190_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[22]~195_combout ))))

	.dataa(\rfif.rdat2[22]~190_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[22]~197_combout ),
	.datad(\rfif.rdat2[22]~195_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~198_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~198 .lut_mask = 16'hF388;
defparam \rfif.rdat2[22]~198 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N27
dffeas \regs[11][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][22] .is_wysiwyg = "true";
defparam \regs[11][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N26
cycloneive_lcell_comb \rfif.rdat2[22]~202 (
// Equation(s):
// \rfif.rdat2[22]~202_combout  = (\rfif.rdat2[22]~201_combout  & (((\regs[11][22]~q ) # (!Instr_IF_16)))) # (!\rfif.rdat2[22]~201_combout  & (\regs[9][22]~q  & ((Instr_IF_16))))

	.dataa(\rfif.rdat2[22]~201_combout ),
	.datab(\regs[9][22]~q ),
	.datac(\regs[11][22]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~202_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~202 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[22]~202 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[22]~203 (
// Equation(s):
// \rfif.rdat2[22]~203_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][22]~q )) # (!Instr_IF_17 & ((\regs[0][22]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[2][22]~q ),
	.datac(\regs[0][22]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~203_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~203 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[22]~203 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[22]~204 (
// Equation(s):
// \rfif.rdat2[22]~204_combout  = (\rfif.rdat2[22]~203_combout  & (((\regs[3][22]~q ) # (!Instr_IF_16)))) # (!\rfif.rdat2[22]~203_combout  & (\regs[1][22]~q  & ((Instr_IF_16))))

	.dataa(\regs[1][22]~q ),
	.datab(\regs[3][22]~q ),
	.datac(\rfif.rdat2[22]~203_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~204_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~204 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[22]~204 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[22]~205 (
// Equation(s):
// \rfif.rdat2[22]~205_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\rfif.rdat2[22]~202_combout )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\rfif.rdat2[22]~204_combout ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[22]~202_combout ),
	.datad(\rfif.rdat2[22]~204_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~205_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~205 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[22]~205 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \rfif.rdat2[22]~200 (
// Equation(s):
// \rfif.rdat2[22]~200_combout  = (\rfif.rdat2[22]~199_combout  & (((\regs[7][22]~q )) # (!Instr_IF_17))) # (!\rfif.rdat2[22]~199_combout  & (Instr_IF_17 & (\regs[6][22]~q )))

	.dataa(\rfif.rdat2[22]~199_combout ),
	.datab(Instr_IF_17),
	.datac(\regs[6][22]~q ),
	.datad(\regs[7][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~200_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~200 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[22]~200 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \rfif.rdat2[22]~207 (
// Equation(s):
// \rfif.rdat2[22]~207_combout  = (\rfif.rdat2[22]~206_combout  & (((\regs[15][22]~q )) # (!Instr_IF_17))) # (!\rfif.rdat2[22]~206_combout  & (Instr_IF_17 & ((\regs[14][22]~q ))))

	.dataa(\rfif.rdat2[22]~206_combout ),
	.datab(Instr_IF_17),
	.datac(\regs[15][22]~q ),
	.datad(\regs[14][22]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~207_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~207 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[22]~207 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \rfif.rdat2[22]~208 (
// Equation(s):
// \rfif.rdat2[22]~208_combout  = (Instr_IF_18 & ((\rfif.rdat2[22]~205_combout  & ((\rfif.rdat2[22]~207_combout ))) # (!\rfif.rdat2[22]~205_combout  & (\rfif.rdat2[22]~200_combout )))) # (!Instr_IF_18 & (\rfif.rdat2[22]~205_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[22]~205_combout ),
	.datac(\rfif.rdat2[22]~200_combout ),
	.datad(\rfif.rdat2[22]~207_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[22]~208_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[22]~208 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[22]~208 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N29
dffeas \regs[20][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][21] .is_wysiwyg = "true";
defparam \regs[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \regs[28][21]~feeder (
// Equation(s):
// \regs[28][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b9),
	.cin(gnd),
	.combout(\regs[28][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N19
dffeas \regs[28][21] (
	.clk(!CLK),
	.d(\regs[28][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][21] .is_wysiwyg = "true";
defparam \regs[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[21]~205 (
// Equation(s):
// \rfif.rdat1[21]~205_combout  = (\rfif.rdat1[21]~204_combout  & (((\regs[28][21]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[21]~204_combout  & (Instr_IF_23 & (\regs[20][21]~q )))

	.dataa(\rfif.rdat1[21]~204_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[20][21]~q ),
	.datad(\regs[28][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~205_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~205 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[21]~205 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N5
dffeas \regs[25][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][21] .is_wysiwyg = "true";
defparam \regs[25][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N9
dffeas \regs[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][21] .is_wysiwyg = "true";
defparam \regs[21][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \rfif.rdat1[21]~202 (
// Equation(s):
// \rfif.rdat1[21]~202_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][21]~q ))) # (!Instr_IF_23 & (\regs[17][21]~q ))))

	.dataa(\regs[17][21]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[21][21]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~202_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~202 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[21]~202 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[21]~203 (
// Equation(s):
// \rfif.rdat1[21]~203_combout  = (Instr_IF_24 & ((\rfif.rdat1[21]~202_combout  & (\regs[29][21]~q )) # (!\rfif.rdat1[21]~202_combout  & ((\regs[25][21]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[21]~202_combout ))))

	.dataa(\regs[29][21]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[25][21]~q ),
	.datad(\rfif.rdat1[21]~202_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~203_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~203 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[21]~203 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[21]~206 (
// Equation(s):
// \rfif.rdat1[21]~206_combout  = (Instr_IF_21 & (((\rfif.rdat1[21]~203_combout ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\rfif.rdat1[21]~205_combout  & ((!Instr_IF_22))))

	.dataa(\rfif.rdat1[21]~205_combout ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[21]~203_combout ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~206_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~206 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[21]~206 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N16
cycloneive_lcell_comb \regs[27][21]~feeder (
// Equation(s):
// \regs[27][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b9),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N17
dffeas \regs[27][21] (
	.clk(!CLK),
	.d(\regs[27][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][21] .is_wysiwyg = "true";
defparam \regs[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N19
dffeas \regs[19][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][21] .is_wysiwyg = "true";
defparam \regs[19][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N17
dffeas \regs[23][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][21] .is_wysiwyg = "true";
defparam \regs[23][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N16
cycloneive_lcell_comb \rfif.rdat1[21]~207 (
// Equation(s):
// \rfif.rdat1[21]~207_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][21]~q ))) # (!Instr_IF_23 & (\regs[19][21]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[19][21]~q ),
	.datac(\regs[23][21]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~207_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~207 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[21]~207 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N7
dffeas \regs[31][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][21] .is_wysiwyg = "true";
defparam \regs[31][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[21]~208 (
// Equation(s):
// \rfif.rdat1[21]~208_combout  = (\rfif.rdat1[21]~207_combout  & (((\regs[31][21]~q ) # (!Instr_IF_24)))) # (!\rfif.rdat1[21]~207_combout  & (\regs[27][21]~q  & (Instr_IF_24)))

	.dataa(\regs[27][21]~q ),
	.datab(\rfif.rdat1[21]~207_combout ),
	.datac(Instr_IF_24),
	.datad(\regs[31][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~208_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~208 .lut_mask = 16'hEC2C;
defparam \rfif.rdat1[21]~208 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N17
dffeas \regs[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][21] .is_wysiwyg = "true";
defparam \regs[22][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas \regs[30][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][21] .is_wysiwyg = "true";
defparam \regs[30][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N11
dffeas \regs[26][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][21] .is_wysiwyg = "true";
defparam \regs[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N19
dffeas \regs[18][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][21] .is_wysiwyg = "true";
defparam \regs[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \rfif.rdat1[21]~200 (
// Equation(s):
// \rfif.rdat1[21]~200_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][21]~q )) # (!Instr_IF_24 & ((\regs[18][21]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][21]~q ),
	.datad(\regs[18][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~200_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~200 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[21]~200 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \rfif.rdat1[21]~201 (
// Equation(s):
// \rfif.rdat1[21]~201_combout  = (Instr_IF_23 & ((\rfif.rdat1[21]~200_combout  & ((\regs[30][21]~q ))) # (!\rfif.rdat1[21]~200_combout  & (\regs[22][21]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[21]~200_combout ))))

	.dataa(\regs[22][21]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[30][21]~q ),
	.datad(\rfif.rdat1[21]~200_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~201_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~201 .lut_mask = 16'hF388;
defparam \rfif.rdat1[21]~201 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \regs[7][21]~feeder (
// Equation(s):
// \regs[7][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b9),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[7][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[7][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N19
dffeas \regs[7][21] (
	.clk(!CLK),
	.d(\regs[7][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][21] .is_wysiwyg = "true";
defparam \regs[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N21
dffeas \regs[6][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][21] .is_wysiwyg = "true";
defparam \regs[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N7
dffeas \regs[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][21] .is_wysiwyg = "true";
defparam \regs[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[21]~212 (
// Equation(s):
// \rfif.rdat1[21]~212_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[6][21]~q )) # (!Instr_IF_22 & ((\regs[4][21]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[6][21]~q ),
	.datad(\regs[4][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~212_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~212 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[21]~212 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \regs[5][21]~feeder (
// Equation(s):
// \regs[5][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b9),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[5][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][21]~feeder .lut_mask = 16'hF0F0;
defparam \regs[5][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N1
dffeas \regs[5][21] (
	.clk(!CLK),
	.d(\regs[5][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][21] .is_wysiwyg = "true";
defparam \regs[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \rfif.rdat1[21]~213 (
// Equation(s):
// \rfif.rdat1[21]~213_combout  = (Instr_IF_21 & ((\rfif.rdat1[21]~212_combout  & (\regs[7][21]~q )) # (!\rfif.rdat1[21]~212_combout  & ((\regs[5][21]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[21]~212_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[7][21]~q ),
	.datac(\rfif.rdat1[21]~212_combout ),
	.datad(\regs[5][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~213_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~213 .lut_mask = 16'hDAD0;
defparam \rfif.rdat1[21]~213 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \regs[3][21]~feeder (
// Equation(s):
// \regs[3][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b9),
	.cin(gnd),
	.combout(\regs[3][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N9
dffeas \regs[3][21] (
	.clk(!CLK),
	.d(\regs[3][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][21] .is_wysiwyg = "true";
defparam \regs[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N31
dffeas \regs[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][21] .is_wysiwyg = "true";
defparam \regs[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[21]~215 (
// Equation(s):
// \rfif.rdat1[21]~215_combout  = (\rfif.rdat1[21]~214_combout  & (((\regs[3][21]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[21]~214_combout  & (Instr_IF_22 & ((\regs[2][21]~q ))))

	.dataa(\rfif.rdat1[21]~214_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[3][21]~q ),
	.datad(\regs[2][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~215_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~215 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[21]~215 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \rfif.rdat1[21]~216 (
// Equation(s):
// \rfif.rdat1[21]~216_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\rfif.rdat1[21]~213_combout )) # (!Instr_IF_23 & ((\rfif.rdat1[21]~215_combout )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[21]~213_combout ),
	.datad(\rfif.rdat1[21]~215_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~216_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~216 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[21]~216 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N27
dffeas \regs[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][21] .is_wysiwyg = "true";
defparam \regs[8][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N13
dffeas \regs[9][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][21] .is_wysiwyg = "true";
defparam \regs[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \rfif.rdat1[21]~210 (
// Equation(s):
// \rfif.rdat1[21]~210_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[9][21]~q ))) # (!Instr_IF_21 & (\regs[8][21]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[8][21]~q ),
	.datad(\regs[9][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~210_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~210 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[21]~210 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N15
dffeas \regs[11][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][21] .is_wysiwyg = "true";
defparam \regs[11][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N5
dffeas \regs[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][21] .is_wysiwyg = "true";
defparam \regs[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[21]~211 (
// Equation(s):
// \rfif.rdat1[21]~211_combout  = (\rfif.rdat1[21]~210_combout  & ((\regs[11][21]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[21]~210_combout  & (((\regs[10][21]~q  & Instr_IF_22))))

	.dataa(\rfif.rdat1[21]~210_combout ),
	.datab(\regs[11][21]~q ),
	.datac(\regs[10][21]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~211_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~211 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[21]~211 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \regs[15][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][21] .is_wysiwyg = "true";
defparam \regs[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N19
dffeas \regs[14][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][21] .is_wysiwyg = "true";
defparam \regs[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N29
dffeas \regs[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][21] .is_wysiwyg = "true";
defparam \regs[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \rfif.rdat1[21]~217 (
// Equation(s):
// \rfif.rdat1[21]~217_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][21]~q )) # (!Instr_IF_22 & ((\regs[12][21]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[14][21]~q ),
	.datad(\regs[12][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~217_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~217 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[21]~217 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N23
dffeas \regs[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][21] .is_wysiwyg = "true";
defparam \regs[13][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \rfif.rdat1[21]~218 (
// Equation(s):
// \rfif.rdat1[21]~218_combout  = (Instr_IF_21 & ((\rfif.rdat1[21]~217_combout  & (\regs[15][21]~q )) # (!\rfif.rdat1[21]~217_combout  & ((\regs[13][21]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[21]~217_combout ))))

	.dataa(\regs[15][21]~q ),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[21]~217_combout ),
	.datad(\regs[13][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[21]~218_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[21]~218 .lut_mask = 16'hBCB0;
defparam \rfif.rdat1[21]~218 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \rfif.rdat2[21]~227 (
// Equation(s):
// \rfif.rdat2[21]~227_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][21]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][21]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][21]~q ),
	.datad(\regs[14][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~227_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~227 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[21]~227 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \rfif.rdat2[21]~228 (
// Equation(s):
// \rfif.rdat2[21]~228_combout  = (Instr_IF_16 & ((\rfif.rdat2[21]~227_combout  & (\regs[15][21]~q )) # (!\rfif.rdat2[21]~227_combout  & ((\regs[13][21]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[21]~227_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[15][21]~q ),
	.datac(\regs[13][21]~q ),
	.datad(\rfif.rdat2[21]~227_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~228_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~228 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[21]~228 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \rfif.rdat2[21]~221 (
// Equation(s):
// \rfif.rdat2[21]~221_combout  = (\rfif.rdat2[21]~220_combout  & (((\regs[11][21]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[21]~220_combout  & (\regs[10][21]~q  & ((Instr_IF_17))))

	.dataa(\rfif.rdat2[21]~220_combout ),
	.datab(\regs[10][21]~q ),
	.datac(\regs[11][21]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~221_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~221 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[21]~221 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \regs[1][21]~feeder (
// Equation(s):
// \regs[1][21]~feeder_combout  = \input_b~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b9),
	.cin(gnd),
	.combout(\regs[1][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][21]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N1
dffeas \regs[1][21] (
	.clk(!CLK),
	.d(\regs[1][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][21] .is_wysiwyg = "true";
defparam \regs[1][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N25
dffeas \regs[0][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][21] .is_wysiwyg = "true";
defparam \regs[0][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \rfif.rdat2[21]~224 (
// Equation(s):
// \rfif.rdat2[21]~224_combout  = (Instr_IF_16 & ((\regs[1][21]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[0][21]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][21]~q ),
	.datac(\regs[0][21]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~224_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~224 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[21]~224 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[21]~225 (
// Equation(s):
// \rfif.rdat2[21]~225_combout  = (Instr_IF_17 & ((\rfif.rdat2[21]~224_combout  & (\regs[3][21]~q )) # (!\rfif.rdat2[21]~224_combout  & ((\regs[2][21]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[21]~224_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[3][21]~q ),
	.datac(\regs[2][21]~q ),
	.datad(\rfif.rdat2[21]~224_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~225_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~225 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[21]~225 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \rfif.rdat2[21]~226 (
// Equation(s):
// \rfif.rdat2[21]~226_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\rfif.rdat2[21]~223_combout )) # (!Instr_IF_18 & ((\rfif.rdat2[21]~225_combout )))))

	.dataa(\rfif.rdat2[21]~223_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[21]~225_combout ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~226_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~226 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[21]~226 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \rfif.rdat2[21]~229 (
// Equation(s):
// \rfif.rdat2[21]~229_combout  = (Instr_IF_19 & ((\rfif.rdat2[21]~226_combout  & (\rfif.rdat2[21]~228_combout )) # (!\rfif.rdat2[21]~226_combout  & ((\rfif.rdat2[21]~221_combout ))))) # (!Instr_IF_19 & (((\rfif.rdat2[21]~226_combout ))))

	.dataa(\rfif.rdat2[21]~228_combout ),
	.datab(\rfif.rdat2[21]~221_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[21]~226_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~229_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~229 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[21]~229 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[21]~217 (
// Equation(s):
// \rfif.rdat2[21]~217_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[23][21]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[19][21]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][21]~q ),
	.datad(\regs[23][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~217_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~217 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[21]~217 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N6
cycloneive_lcell_comb \rfif.rdat2[21]~218 (
// Equation(s):
// \rfif.rdat2[21]~218_combout  = (\rfif.rdat2[21]~217_combout  & (((\regs[31][21]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[21]~217_combout  & (\regs[27][21]~q  & ((Instr_IF_19))))

	.dataa(\regs[27][21]~q ),
	.datab(\rfif.rdat2[21]~217_combout ),
	.datac(\regs[31][21]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~218_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~218 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[21]~218 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \rfif.rdat2[21]~210 (
// Equation(s):
// \rfif.rdat2[21]~210_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][21]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][21]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][21]~q ),
	.datad(\regs[26][21]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~210_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~210 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[21]~210 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \rfif.rdat2[21]~211 (
// Equation(s):
// \rfif.rdat2[21]~211_combout  = (Instr_IF_18 & ((\rfif.rdat2[21]~210_combout  & (\regs[30][21]~q )) # (!\rfif.rdat2[21]~210_combout  & ((\regs[22][21]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[21]~210_combout ))))

	.dataa(\regs[30][21]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][21]~q ),
	.datad(\rfif.rdat2[21]~210_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~211_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~211 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[21]~211 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas \regs[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][21] .is_wysiwyg = "true";
defparam \regs[29][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N11
dffeas \regs[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][21] .is_wysiwyg = "true";
defparam \regs[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[21]~212 (
// Equation(s):
// \rfif.rdat2[21]~212_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[21][21]~q )) # (!Instr_IF_18 & ((\regs[17][21]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[21][21]~q ),
	.datac(\regs[17][21]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~212_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~212 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[21]~212 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[21]~213 (
// Equation(s):
// \rfif.rdat2[21]~213_combout  = (Instr_IF_19 & ((\rfif.rdat2[21]~212_combout  & ((\regs[29][21]~q ))) # (!\rfif.rdat2[21]~212_combout  & (\regs[25][21]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[21]~212_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][21]~q ),
	.datac(\regs[29][21]~q ),
	.datad(\rfif.rdat2[21]~212_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~213_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~213 .lut_mask = 16'hF588;
defparam \rfif.rdat2[21]~213 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \rfif.rdat2[21]~216 (
// Equation(s):
// \rfif.rdat2[21]~216_combout  = (Instr_IF_16 & (((Instr_IF_17) # (\rfif.rdat2[21]~213_combout )))) # (!Instr_IF_16 & (\rfif.rdat2[21]~215_combout  & (!Instr_IF_17)))

	.dataa(\rfif.rdat2[21]~215_combout ),
	.datab(Instr_IF_16),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[21]~213_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~216_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~216 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[21]~216 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \rfif.rdat2[21]~219 (
// Equation(s):
// \rfif.rdat2[21]~219_combout  = (Instr_IF_17 & ((\rfif.rdat2[21]~216_combout  & (\rfif.rdat2[21]~218_combout )) # (!\rfif.rdat2[21]~216_combout  & ((\rfif.rdat2[21]~211_combout ))))) # (!Instr_IF_17 & (((\rfif.rdat2[21]~216_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[21]~218_combout ),
	.datac(\rfif.rdat2[21]~211_combout ),
	.datad(\rfif.rdat2[21]~216_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[21]~219_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[21]~219 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[21]~219 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N17
dffeas \regs[27][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][20] .is_wysiwyg = "true";
defparam \regs[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N13
dffeas \regs[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][20] .is_wysiwyg = "true";
defparam \regs[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[20]~227 (
// Equation(s):
// \rfif.rdat1[20]~227_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][20]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][20]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][20]~q ),
	.datad(\regs[19][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~227_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~227 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[20]~227 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N27
dffeas \regs[23][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][20] .is_wysiwyg = "true";
defparam \regs[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N25
dffeas \regs[31][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][20] .is_wysiwyg = "true";
defparam \regs[31][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N26
cycloneive_lcell_comb \rfif.rdat1[20]~228 (
// Equation(s):
// \rfif.rdat1[20]~228_combout  = (Instr_IF_23 & ((\rfif.rdat1[20]~227_combout  & ((\regs[31][20]~q ))) # (!\rfif.rdat1[20]~227_combout  & (\regs[23][20]~q )))) # (!Instr_IF_23 & (\rfif.rdat1[20]~227_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[20]~227_combout ),
	.datac(\regs[23][20]~q ),
	.datad(\regs[31][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~228_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~228 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[20]~228 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N21
dffeas \regs[21][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][20] .is_wysiwyg = "true";
defparam \regs[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N15
dffeas \regs[29][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][20] .is_wysiwyg = "true";
defparam \regs[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N3
dffeas \regs[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][20] .is_wysiwyg = "true";
defparam \regs[17][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \regs[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][20] .is_wysiwyg = "true";
defparam \regs[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[20]~220 (
// Equation(s):
// \rfif.rdat1[20]~220_combout  = (Instr_IF_24 & (((\regs[25][20]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][20]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][20]~q ),
	.datac(\regs[25][20]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~220_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~220 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[20]~220 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[20]~221 (
// Equation(s):
// \rfif.rdat1[20]~221_combout  = (Instr_IF_23 & ((\rfif.rdat1[20]~220_combout  & ((\regs[29][20]~q ))) # (!\rfif.rdat1[20]~220_combout  & (\regs[21][20]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[20]~220_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[21][20]~q ),
	.datac(\regs[29][20]~q ),
	.datad(\rfif.rdat1[20]~220_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~221_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~221 .lut_mask = 16'hF588;
defparam \rfif.rdat1[20]~221 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \regs[24][20]~feeder (
// Equation(s):
// \regs[24][20]~feeder_combout  = \input_b~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \regs[24][20] (
	.clk(!CLK),
	.d(\regs[24][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][20] .is_wysiwyg = "true";
defparam \regs[24][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N9
dffeas \regs[20][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][20] .is_wysiwyg = "true";
defparam \regs[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[20]~224 (
// Equation(s):
// \rfif.rdat1[20]~224_combout  = (Instr_IF_23 & (((\regs[20][20]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][20]~q  & ((!Instr_IF_24))))

	.dataa(\regs[16][20]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][20]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~224_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~224 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[20]~224 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \rfif.rdat1[20]~225 (
// Equation(s):
// \rfif.rdat1[20]~225_combout  = (\rfif.rdat1[20]~224_combout  & ((\regs[28][20]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[20]~224_combout  & (((\regs[24][20]~q  & Instr_IF_24))))

	.dataa(\regs[28][20]~q ),
	.datab(\regs[24][20]~q ),
	.datac(\rfif.rdat1[20]~224_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~225_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~225 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[20]~225 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \regs[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][20] .is_wysiwyg = "true";
defparam \regs[18][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N13
dffeas \regs[22][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][20] .is_wysiwyg = "true";
defparam \regs[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \rfif.rdat1[20]~222 (
// Equation(s):
// \rfif.rdat1[20]~222_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][20]~q ))) # (!Instr_IF_23 & (\regs[18][20]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[18][20]~q ),
	.datac(\regs[22][20]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~222_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~222 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[20]~222 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N9
dffeas \regs[26][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][20] .is_wysiwyg = "true";
defparam \regs[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N3
dffeas \regs[30][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][20] .is_wysiwyg = "true";
defparam \regs[30][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[20]~223 (
// Equation(s):
// \rfif.rdat1[20]~223_combout  = (Instr_IF_24 & ((\rfif.rdat1[20]~222_combout  & ((\regs[30][20]~q ))) # (!\rfif.rdat1[20]~222_combout  & (\regs[26][20]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[20]~222_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[20]~222_combout ),
	.datac(\regs[26][20]~q ),
	.datad(\regs[30][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~223_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~223 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[20]~223 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \rfif.rdat1[20]~226 (
// Equation(s):
// \rfif.rdat1[20]~226_combout  = (Instr_IF_22 & (((\rfif.rdat1[20]~223_combout ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\rfif.rdat1[20]~225_combout  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[20]~225_combout ),
	.datac(\rfif.rdat1[20]~223_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~226_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~226 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[20]~226 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N25
dffeas \regs[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][20] .is_wysiwyg = "true";
defparam \regs[10][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N23
dffeas \regs[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][20] .is_wysiwyg = "true";
defparam \regs[8][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[20]~232 (
// Equation(s):
// \rfif.rdat1[20]~232_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][20]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][20]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][20]~q ),
	.datad(\regs[8][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~232_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~232 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[20]~232 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N1
dffeas \regs[9][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][20] .is_wysiwyg = "true";
defparam \regs[9][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[20]~233 (
// Equation(s):
// \rfif.rdat1[20]~233_combout  = (\rfif.rdat1[20]~232_combout  & ((\regs[11][20]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[20]~232_combout  & (((\regs[9][20]~q  & Instr_IF_21))))

	.dataa(\regs[11][20]~q ),
	.datab(\rfif.rdat1[20]~232_combout ),
	.datac(\regs[9][20]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~233_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~233 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[20]~233 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N19
dffeas \regs[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][20] .is_wysiwyg = "true";
defparam \regs[3][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N5
dffeas \regs[1][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][20] .is_wysiwyg = "true";
defparam \regs[1][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N21
dffeas \regs[0][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][20] .is_wysiwyg = "true";
defparam \regs[0][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \regs[2][20]~feeder (
// Equation(s):
// \regs[2][20]~feeder_combout  = \input_b~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N7
dffeas \regs[2][20] (
	.clk(!CLK),
	.d(\regs[2][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][20] .is_wysiwyg = "true";
defparam \regs[2][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[20]~234 (
// Equation(s):
// \rfif.rdat1[20]~234_combout  = (Instr_IF_22 & (((Instr_IF_21) # (\regs[2][20]~q )))) # (!Instr_IF_22 & (\regs[0][20]~q  & (!Instr_IF_21)))

	.dataa(Instr_IF_22),
	.datab(\regs[0][20]~q ),
	.datac(Instr_IF_21),
	.datad(\regs[2][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~234_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~234 .lut_mask = 16'hAEA4;
defparam \rfif.rdat1[20]~234 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[20]~235 (
// Equation(s):
// \rfif.rdat1[20]~235_combout  = (Instr_IF_21 & ((\rfif.rdat1[20]~234_combout  & (\regs[3][20]~q )) # (!\rfif.rdat1[20]~234_combout  & ((\regs[1][20]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[20]~234_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[3][20]~q ),
	.datac(\regs[1][20]~q ),
	.datad(\rfif.rdat1[20]~234_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~235_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~235 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[20]~235 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \rfif.rdat1[20]~236 (
// Equation(s):
// \rfif.rdat1[20]~236_combout  = (Instr_IF_24 & ((\rfif.rdat1[20]~233_combout ) # ((Instr_IF_23)))) # (!Instr_IF_24 & (((!Instr_IF_23 & \rfif.rdat1[20]~235_combout ))))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[20]~233_combout ),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[20]~235_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~236_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~236 .lut_mask = 16'hADA8;
defparam \rfif.rdat1[20]~236 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N15
dffeas \regs[15][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][20] .is_wysiwyg = "true";
defparam \regs[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N7
dffeas \regs[13][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][20] .is_wysiwyg = "true";
defparam \regs[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \rfif.rdat1[20]~237 (
// Equation(s):
// \rfif.rdat1[20]~237_combout  = (Instr_IF_21 & (((\regs[13][20]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][20]~q  & ((!Instr_IF_22))))

	.dataa(\regs[12][20]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][20]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~237_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~237 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[20]~237 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \regs[14][20]~feeder (
// Equation(s):
// \regs[14][20]~feeder_combout  = \input_b~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N17
dffeas \regs[14][20] (
	.clk(!CLK),
	.d(\regs[14][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][20] .is_wysiwyg = "true";
defparam \regs[14][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \rfif.rdat1[20]~238 (
// Equation(s):
// \rfif.rdat1[20]~238_combout  = (\rfif.rdat1[20]~237_combout  & ((\regs[15][20]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[20]~237_combout  & (((Instr_IF_22 & \regs[14][20]~q ))))

	.dataa(\regs[15][20]~q ),
	.datab(\rfif.rdat1[20]~237_combout ),
	.datac(Instr_IF_22),
	.datad(\regs[14][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~238_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~238 .lut_mask = 16'hBC8C;
defparam \rfif.rdat1[20]~238 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \regs[6][20]~feeder (
// Equation(s):
// \regs[6][20]~feeder_combout  = \input_b~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][20]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N11
dffeas \regs[6][20] (
	.clk(!CLK),
	.d(\regs[6][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][20] .is_wysiwyg = "true";
defparam \regs[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N1
dffeas \regs[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][20] .is_wysiwyg = "true";
defparam \regs[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N23
dffeas \regs[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][20] .is_wysiwyg = "true";
defparam \regs[5][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \rfif.rdat1[20]~230 (
// Equation(s):
// \rfif.rdat1[20]~230_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][20]~q ))) # (!Instr_IF_21 & (\regs[4][20]~q ))))

	.dataa(\regs[4][20]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][20]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~230_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~230 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[20]~230 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \rfif.rdat1[20]~231 (
// Equation(s):
// \rfif.rdat1[20]~231_combout  = (Instr_IF_22 & ((\rfif.rdat1[20]~230_combout  & ((\regs[7][20]~q ))) # (!\rfif.rdat1[20]~230_combout  & (\regs[6][20]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[20]~230_combout ))))

	.dataa(\regs[6][20]~q ),
	.datab(\regs[7][20]~q ),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[20]~230_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[20]~231_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[20]~231 .lut_mask = 16'hCFA0;
defparam \rfif.rdat1[20]~231 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[20]~238 (
// Equation(s):
// \rfif.rdat2[20]~238_combout  = (Instr_IF_19 & ((\regs[27][20]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[19][20]~q  & !Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][20]~q ),
	.datac(\regs[19][20]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~238_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~238 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[20]~238 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \rfif.rdat2[20]~239 (
// Equation(s):
// \rfif.rdat2[20]~239_combout  = (Instr_IF_18 & ((\rfif.rdat2[20]~238_combout  & ((\regs[31][20]~q ))) # (!\rfif.rdat2[20]~238_combout  & (\regs[23][20]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[20]~238_combout ))))

	.dataa(\regs[23][20]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[31][20]~q ),
	.datad(\rfif.rdat2[20]~238_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~239_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~239 .lut_mask = 16'hF388;
defparam \rfif.rdat2[20]~239 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[20]~233 (
// Equation(s):
// \rfif.rdat2[20]~233_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][20]~q ))) # (!Instr_IF_18 & (\regs[18][20]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][20]~q ),
	.datad(\regs[22][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~233_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~233 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[20]~233 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \rfif.rdat2[20]~234 (
// Equation(s):
// \rfif.rdat2[20]~234_combout  = (\rfif.rdat2[20]~233_combout  & (((\regs[30][20]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[20]~233_combout  & (\regs[26][20]~q  & ((Instr_IF_19))))

	.dataa(\regs[26][20]~q ),
	.datab(\rfif.rdat2[20]~233_combout ),
	.datac(\regs[30][20]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~234_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~234 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[20]~234 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N13
dffeas \regs[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][20] .is_wysiwyg = "true";
defparam \regs[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \rfif.rdat2[20]~236 (
// Equation(s):
// \rfif.rdat2[20]~236_combout  = (\rfif.rdat2[20]~235_combout  & (((\regs[28][20]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[20]~235_combout  & (\regs[24][20]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[20]~235_combout ),
	.datab(\regs[24][20]~q ),
	.datac(\regs[28][20]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~236_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~236 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[20]~236 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \rfif.rdat2[20]~237 (
// Equation(s):
// \rfif.rdat2[20]~237_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\rfif.rdat2[20]~234_combout )))) # (!Instr_IF_17 & (!Instr_IF_16 & ((\rfif.rdat2[20]~236_combout ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[20]~234_combout ),
	.datad(\rfif.rdat2[20]~236_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~237_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~237 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[20]~237 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[20]~231 (
// Equation(s):
// \rfif.rdat2[20]~231_combout  = (Instr_IF_19 & ((\regs[25][20]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\regs[17][20]~q  & !Instr_IF_18))))

	.dataa(\regs[25][20]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[17][20]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~231_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~231 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[20]~231 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \rfif.rdat2[20]~232 (
// Equation(s):
// \rfif.rdat2[20]~232_combout  = (\rfif.rdat2[20]~231_combout  & ((\regs[29][20]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[20]~231_combout  & (((\regs[21][20]~q  & Instr_IF_18))))

	.dataa(\regs[29][20]~q ),
	.datab(\rfif.rdat2[20]~231_combout ),
	.datac(\regs[21][20]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~232_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~232 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[20]~232 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \rfif.rdat2[20]~240 (
// Equation(s):
// \rfif.rdat2[20]~240_combout  = (\rfif.rdat2[20]~237_combout  & ((\rfif.rdat2[20]~239_combout ) # ((!Instr_IF_16)))) # (!\rfif.rdat2[20]~237_combout  & (((\rfif.rdat2[20]~232_combout  & Instr_IF_16))))

	.dataa(\rfif.rdat2[20]~239_combout ),
	.datab(\rfif.rdat2[20]~237_combout ),
	.datac(\rfif.rdat2[20]~232_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~240_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~240 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[20]~240 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[20]~245 (
// Equation(s):
// \rfif.rdat2[20]~245_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][20]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][20]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][20]~q ),
	.datad(\regs[2][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~245_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~245 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[20]~245 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[20]~246 (
// Equation(s):
// \rfif.rdat2[20]~246_combout  = (Instr_IF_16 & ((\rfif.rdat2[20]~245_combout  & ((\regs[3][20]~q ))) # (!\rfif.rdat2[20]~245_combout  & (\regs[1][20]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[20]~245_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][20]~q ),
	.datac(\regs[3][20]~q ),
	.datad(\rfif.rdat2[20]~245_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~246_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~246 .lut_mask = 16'hF588;
defparam \rfif.rdat2[20]~246 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[20]~243 (
// Equation(s):
// \rfif.rdat2[20]~243_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][20]~q ))) # (!Instr_IF_17 & (\regs[8][20]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][20]~q ),
	.datad(\regs[10][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~243_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~243 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[20]~243 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N31
dffeas \regs[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][20] .is_wysiwyg = "true";
defparam \regs[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[20]~244 (
// Equation(s):
// \rfif.rdat2[20]~244_combout  = (Instr_IF_16 & ((\rfif.rdat2[20]~243_combout  & (\regs[11][20]~q )) # (!\rfif.rdat2[20]~243_combout  & ((\regs[9][20]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[20]~243_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[20]~243_combout ),
	.datac(\regs[11][20]~q ),
	.datad(\regs[9][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~244_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~244 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[20]~244 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \rfif.rdat2[20]~247 (
// Equation(s):
// \rfif.rdat2[20]~247_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\rfif.rdat2[20]~244_combout ))) # (!Instr_IF_19 & (\rfif.rdat2[20]~246_combout ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[20]~246_combout ),
	.datad(\rfif.rdat2[20]~244_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~247_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~247 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[20]~247 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N17
dffeas \regs[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][20] .is_wysiwyg = "true";
defparam \regs[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \rfif.rdat2[20]~241 (
// Equation(s):
// \rfif.rdat2[20]~241_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][20]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][20]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][20]~q ),
	.datad(\regs[5][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~241_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~241 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[20]~241 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[20]~242 (
// Equation(s):
// \rfif.rdat2[20]~242_combout  = (Instr_IF_17 & ((\rfif.rdat2[20]~241_combout  & ((\regs[7][20]~q ))) # (!\rfif.rdat2[20]~241_combout  & (\regs[6][20]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[20]~241_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[6][20]~q ),
	.datac(\regs[7][20]~q ),
	.datad(\rfif.rdat2[20]~241_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~242_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~242 .lut_mask = 16'hF588;
defparam \rfif.rdat2[20]~242 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \regs[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][20] .is_wysiwyg = "true";
defparam \regs[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \rfif.rdat2[20]~248 (
// Equation(s):
// \rfif.rdat2[20]~248_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[13][20]~q ))) # (!Instr_IF_16 & (\regs[12][20]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][20]~q ),
	.datad(\regs[13][20]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~248_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~248 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[20]~248 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[20]~249 (
// Equation(s):
// \rfif.rdat2[20]~249_combout  = (Instr_IF_17 & ((\rfif.rdat2[20]~248_combout  & (\regs[15][20]~q )) # (!\rfif.rdat2[20]~248_combout  & ((\regs[14][20]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[20]~248_combout ))))

	.dataa(\regs[15][20]~q ),
	.datab(\regs[14][20]~q ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[20]~248_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~249_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~249 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[20]~249 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[20]~250 (
// Equation(s):
// \rfif.rdat2[20]~250_combout  = (\rfif.rdat2[20]~247_combout  & (((\rfif.rdat2[20]~249_combout ) # (!Instr_IF_18)))) # (!\rfif.rdat2[20]~247_combout  & (\rfif.rdat2[20]~242_combout  & (Instr_IF_18)))

	.dataa(\rfif.rdat2[20]~247_combout ),
	.datab(\rfif.rdat2[20]~242_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[20]~249_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[20]~250_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[20]~250 .lut_mask = 16'hEA4A;
defparam \rfif.rdat2[20]~250 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \regs[26][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][19] .is_wysiwyg = "true";
defparam \regs[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N31
dffeas \regs[18][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][19] .is_wysiwyg = "true";
defparam \regs[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \rfif.rdat1[19]~240 (
// Equation(s):
// \rfif.rdat1[19]~240_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][19]~q )) # (!Instr_IF_24 & ((\regs[18][19]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][19]~q ),
	.datad(\regs[18][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~240_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~240 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[19]~240 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N1
dffeas \regs[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][19] .is_wysiwyg = "true";
defparam \regs[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \regs[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][19] .is_wysiwyg = "true";
defparam \regs[22][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[19]~241 (
// Equation(s):
// \rfif.rdat1[19]~241_combout  = (Instr_IF_23 & ((\rfif.rdat1[19]~240_combout  & (\regs[30][19]~q )) # (!\rfif.rdat1[19]~240_combout  & ((\regs[22][19]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[19]~240_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[19]~240_combout ),
	.datac(\regs[30][19]~q ),
	.datad(\regs[22][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~241_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~241 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[19]~241 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N23
dffeas \regs[19][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][19] .is_wysiwyg = "true";
defparam \regs[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \regs[23][19]~feeder (
// Equation(s):
// \regs[23][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[23][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[23][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N17
dffeas \regs[23][19] (
	.clk(!CLK),
	.d(\regs[23][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][19] .is_wysiwyg = "true";
defparam \regs[23][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[19]~247 (
// Equation(s):
// \rfif.rdat1[19]~247_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][19]~q ))) # (!Instr_IF_23 & (\regs[19][19]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[19][19]~q ),
	.datad(\regs[23][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~247_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~247 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[19]~247 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N15
dffeas \regs[27][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][19] .is_wysiwyg = "true";
defparam \regs[27][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N13
dffeas \regs[31][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][19] .is_wysiwyg = "true";
defparam \regs[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[19]~248 (
// Equation(s):
// \rfif.rdat1[19]~248_combout  = (Instr_IF_24 & ((\rfif.rdat1[19]~247_combout  & ((\regs[31][19]~q ))) # (!\rfif.rdat1[19]~247_combout  & (\regs[27][19]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[19]~247_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[19]~247_combout ),
	.datac(\regs[27][19]~q ),
	.datad(\regs[31][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~248_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~248 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[19]~248 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N5
dffeas \regs[20][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][19] .is_wysiwyg = "true";
defparam \regs[20][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \regs[28][19]~feeder (
// Equation(s):
// \regs[28][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N27
dffeas \regs[28][19] (
	.clk(!CLK),
	.d(\regs[28][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][19] .is_wysiwyg = "true";
defparam \regs[28][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[19]~245 (
// Equation(s):
// \rfif.rdat1[19]~245_combout  = (\rfif.rdat1[19]~244_combout  & (((\regs[28][19]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[19]~244_combout  & (Instr_IF_23 & (\regs[20][19]~q )))

	.dataa(\rfif.rdat1[19]~244_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[20][19]~q ),
	.datad(\regs[28][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~245_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~245 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[19]~245 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N9
dffeas \regs[25][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][19] .is_wysiwyg = "true";
defparam \regs[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N19
dffeas \regs[29][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][19] .is_wysiwyg = "true";
defparam \regs[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[19]~243 (
// Equation(s):
// \rfif.rdat1[19]~243_combout  = (\rfif.rdat1[19]~242_combout  & (((\regs[29][19]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[19]~242_combout  & (Instr_IF_24 & (\regs[25][19]~q )))

	.dataa(\rfif.rdat1[19]~242_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[25][19]~q ),
	.datad(\regs[29][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~243_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~243 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[19]~243 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[19]~246 (
// Equation(s):
// \rfif.rdat1[19]~246_combout  = (Instr_IF_21 & (((Instr_IF_22) # (\rfif.rdat1[19]~243_combout )))) # (!Instr_IF_21 & (\rfif.rdat1[19]~245_combout  & (!Instr_IF_22)))

	.dataa(\rfif.rdat1[19]~245_combout ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[19]~243_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~246_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~246 .lut_mask = 16'hCEC2;
defparam \rfif.rdat1[19]~246 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \regs[3][19]~feeder (
// Equation(s):
// \regs[3][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b11),
	.cin(gnd),
	.combout(\regs[3][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N5
dffeas \regs[3][19] (
	.clk(!CLK),
	.d(\regs[3][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][19] .is_wysiwyg = "true";
defparam \regs[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \regs[0][19]~feeder (
// Equation(s):
// \regs[0][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b11),
	.cin(gnd),
	.combout(\regs[0][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[0][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[0][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N9
dffeas \regs[0][19] (
	.clk(!CLK),
	.d(\regs[0][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][19] .is_wysiwyg = "true";
defparam \regs[0][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \rfif.rdat1[19]~254 (
// Equation(s):
// \rfif.rdat1[19]~254_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][19]~q )) # (!Instr_IF_21 & ((\regs[0][19]~q )))))

	.dataa(\regs[1][19]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[0][19]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~254_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~254 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[19]~254 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[19]~255 (
// Equation(s):
// \rfif.rdat1[19]~255_combout  = (Instr_IF_22 & ((\rfif.rdat1[19]~254_combout  & ((\regs[3][19]~q ))) # (!\rfif.rdat1[19]~254_combout  & (\regs[2][19]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[19]~254_combout ))))

	.dataa(\regs[2][19]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[3][19]~q ),
	.datad(\rfif.rdat1[19]~254_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~255_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~255 .lut_mask = 16'hF388;
defparam \rfif.rdat1[19]~255 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \regs[5][19]~feeder (
// Equation(s):
// \regs[5][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[5][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[5][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N5
dffeas \regs[5][19] (
	.clk(!CLK),
	.d(\regs[5][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][19] .is_wysiwyg = "true";
defparam \regs[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \regs[7][19]~feeder (
// Equation(s):
// \regs[7][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[7][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[7][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N31
dffeas \regs[7][19] (
	.clk(!CLK),
	.d(\regs[7][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][19] .is_wysiwyg = "true";
defparam \regs[7][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \rfif.rdat1[19]~253 (
// Equation(s):
// \rfif.rdat1[19]~253_combout  = (\rfif.rdat1[19]~252_combout  & (((\regs[7][19]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[19]~252_combout  & (Instr_IF_21 & (\regs[5][19]~q )))

	.dataa(\rfif.rdat1[19]~252_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[5][19]~q ),
	.datad(\regs[7][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~253_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~253 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[19]~253 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \rfif.rdat1[19]~256 (
// Equation(s):
// \rfif.rdat1[19]~256_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\rfif.rdat1[19]~253_combout ))) # (!Instr_IF_23 & (\rfif.rdat1[19]~255_combout ))))

	.dataa(\rfif.rdat1[19]~255_combout ),
	.datab(Instr_IF_24),
	.datac(Instr_IF_23),
	.datad(\rfif.rdat1[19]~253_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~256_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~256 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[19]~256 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \regs[9][19]~feeder (
// Equation(s):
// \regs[9][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b11),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][19]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N21
dffeas \regs[9][19] (
	.clk(!CLK),
	.d(\regs[9][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][19] .is_wysiwyg = "true";
defparam \regs[9][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[19]~250 (
// Equation(s):
// \rfif.rdat1[19]~250_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[9][19]~q ))) # (!Instr_IF_21 & (\regs[8][19]~q ))))

	.dataa(\regs[8][19]~q ),
	.datab(\regs[9][19]~q ),
	.datac(Instr_IF_22),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~250_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~250 .lut_mask = 16'hFC0A;
defparam \rfif.rdat1[19]~250 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N13
dffeas \regs[11][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][19] .is_wysiwyg = "true";
defparam \regs[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N21
dffeas \regs[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][19] .is_wysiwyg = "true";
defparam \regs[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[19]~251 (
// Equation(s):
// \rfif.rdat1[19]~251_combout  = (Instr_IF_22 & ((\rfif.rdat1[19]~250_combout  & (\regs[11][19]~q )) # (!\rfif.rdat1[19]~250_combout  & ((\regs[10][19]~q ))))) # (!Instr_IF_22 & (\rfif.rdat1[19]~250_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[19]~250_combout ),
	.datac(\regs[11][19]~q ),
	.datad(\regs[10][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~251_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~251 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[19]~251 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N25
dffeas \regs[15][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][19] .is_wysiwyg = "true";
defparam \regs[15][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \regs[13][19]~feeder (
// Equation(s):
// \regs[13][19]~feeder_combout  = \input_b~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b11),
	.cin(gnd),
	.combout(\regs[13][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][19]~feeder .lut_mask = 16'hFF00;
defparam \regs[13][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N25
dffeas \regs[13][19] (
	.clk(!CLK),
	.d(\regs[13][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][19] .is_wysiwyg = "true";
defparam \regs[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N1
dffeas \regs[14][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][19] .is_wysiwyg = "true";
defparam \regs[14][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N7
dffeas \regs[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][19] .is_wysiwyg = "true";
defparam \regs[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[19]~257 (
// Equation(s):
// \rfif.rdat1[19]~257_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][19]~q )) # (!Instr_IF_22 & ((\regs[12][19]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[14][19]~q ),
	.datad(\regs[12][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~257_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~257 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[19]~257 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[19]~258 (
// Equation(s):
// \rfif.rdat1[19]~258_combout  = (Instr_IF_21 & ((\rfif.rdat1[19]~257_combout  & (\regs[15][19]~q )) # (!\rfif.rdat1[19]~257_combout  & ((\regs[13][19]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[19]~257_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[15][19]~q ),
	.datac(\regs[13][19]~q ),
	.datad(\rfif.rdat1[19]~257_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[19]~258_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[19]~258 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[19]~258 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[19]~266 (
// Equation(s):
// \rfif.rdat2[19]~266_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[1][19]~q )) # (!Instr_IF_16 & ((\regs[0][19]~q )))))

	.dataa(\regs[1][19]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[0][19]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~266_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~266 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[19]~266 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[19]~267 (
// Equation(s):
// \rfif.rdat2[19]~267_combout  = (Instr_IF_17 & ((\rfif.rdat2[19]~266_combout  & ((\regs[3][19]~q ))) # (!\rfif.rdat2[19]~266_combout  & (\regs[2][19]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[19]~266_combout ))))

	.dataa(\regs[2][19]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[3][19]~q ),
	.datad(\rfif.rdat2[19]~266_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~267_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~267 .lut_mask = 16'hF388;
defparam \rfif.rdat2[19]~267 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N5
dffeas \regs[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][19] .is_wysiwyg = "true";
defparam \regs[4][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N11
dffeas \regs[6][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][19] .is_wysiwyg = "true";
defparam \regs[6][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \rfif.rdat2[19]~264 (
// Equation(s):
// \rfif.rdat2[19]~264_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][19]~q ))) # (!Instr_IF_17 & (\regs[4][19]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][19]~q ),
	.datad(\regs[6][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~264_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~264 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[19]~264 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[19]~265 (
// Equation(s):
// \rfif.rdat2[19]~265_combout  = (Instr_IF_16 & ((\rfif.rdat2[19]~264_combout  & (\regs[7][19]~q )) # (!\rfif.rdat2[19]~264_combout  & ((\regs[5][19]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[19]~264_combout ))))

	.dataa(\regs[7][19]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[5][19]~q ),
	.datad(\rfif.rdat2[19]~264_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~265_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~265 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[19]~265 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[19]~268 (
// Equation(s):
// \rfif.rdat2[19]~268_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\rfif.rdat2[19]~265_combout )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\rfif.rdat2[19]~267_combout )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[19]~267_combout ),
	.datad(\rfif.rdat2[19]~265_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~268_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~268 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[19]~268 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N11
dffeas \regs[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][19] .is_wysiwyg = "true";
defparam \regs[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \rfif.rdat2[19]~262 (
// Equation(s):
// \rfif.rdat2[19]~262_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][19]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][19]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][19]~q ),
	.datad(\regs[9][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~262_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~262 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[19]~262 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \rfif.rdat2[19]~263 (
// Equation(s):
// \rfif.rdat2[19]~263_combout  = (Instr_IF_17 & ((\rfif.rdat2[19]~262_combout  & (\regs[11][19]~q )) # (!\rfif.rdat2[19]~262_combout  & ((\regs[10][19]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[19]~262_combout ))))

	.dataa(\regs[11][19]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[10][19]~q ),
	.datad(\rfif.rdat2[19]~262_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~263_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~263 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[19]~263 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[19]~270 (
// Equation(s):
// \rfif.rdat2[19]~270_combout  = (\rfif.rdat2[19]~269_combout  & (((\regs[15][19]~q ) # (!Instr_IF_16)))) # (!\rfif.rdat2[19]~269_combout  & (\regs[13][19]~q  & ((Instr_IF_16))))

	.dataa(\rfif.rdat2[19]~269_combout ),
	.datab(\regs[13][19]~q ),
	.datac(\regs[15][19]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~270_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~270 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[19]~270 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[19]~271 (
// Equation(s):
// \rfif.rdat2[19]~271_combout  = (\rfif.rdat2[19]~268_combout  & (((\rfif.rdat2[19]~270_combout ) # (!Instr_IF_19)))) # (!\rfif.rdat2[19]~268_combout  & (\rfif.rdat2[19]~263_combout  & (Instr_IF_19)))

	.dataa(\rfif.rdat2[19]~268_combout ),
	.datab(\rfif.rdat2[19]~263_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[19]~270_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~271_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~271 .lut_mask = 16'hEA4A;
defparam \rfif.rdat2[19]~271 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \rfif.rdat2[19]~252 (
// Equation(s):
// \rfif.rdat2[19]~252_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][19]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][19]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][19]~q ),
	.datad(\regs[26][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~252_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~252 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[19]~252 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \rfif.rdat2[19]~253 (
// Equation(s):
// \rfif.rdat2[19]~253_combout  = (Instr_IF_18 & ((\rfif.rdat2[19]~252_combout  & (\regs[30][19]~q )) # (!\rfif.rdat2[19]~252_combout  & ((\regs[22][19]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[19]~252_combout ))))

	.dataa(\regs[30][19]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][19]~q ),
	.datad(\rfif.rdat2[19]~252_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~253_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~253 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[19]~253 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[19]~259 (
// Equation(s):
// \rfif.rdat2[19]~259_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[23][19]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[19][19]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][19]~q ),
	.datad(\regs[23][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~259_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~259 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[19]~259 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[19]~260 (
// Equation(s):
// \rfif.rdat2[19]~260_combout  = (Instr_IF_19 & ((\rfif.rdat2[19]~259_combout  & ((\regs[31][19]~q ))) # (!\rfif.rdat2[19]~259_combout  & (\regs[27][19]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[19]~259_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][19]~q ),
	.datac(\regs[31][19]~q ),
	.datad(\rfif.rdat2[19]~259_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~260_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~260 .lut_mask = 16'hF588;
defparam \rfif.rdat2[19]~260 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas \regs[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][19] .is_wysiwyg = "true";
defparam \regs[17][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N1
dffeas \regs[21][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][19] .is_wysiwyg = "true";
defparam \regs[21][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[19]~254 (
// Equation(s):
// \rfif.rdat2[19]~254_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][19]~q ))) # (!Instr_IF_18 & (\regs[17][19]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][19]~q ),
	.datad(\regs[21][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~254_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~254 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[19]~254 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[19]~255 (
// Equation(s):
// \rfif.rdat2[19]~255_combout  = (Instr_IF_19 & ((\rfif.rdat2[19]~254_combout  & ((\regs[29][19]~q ))) # (!\rfif.rdat2[19]~254_combout  & (\regs[25][19]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[19]~254_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][19]~q ),
	.datac(\regs[29][19]~q ),
	.datad(\rfif.rdat2[19]~254_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~255_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~255 .lut_mask = 16'hF588;
defparam \rfif.rdat2[19]~255 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N21
dffeas \regs[24][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][19] .is_wysiwyg = "true";
defparam \regs[24][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \regs[16][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][19] .is_wysiwyg = "true";
defparam \regs[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[19]~256 (
// Equation(s):
// \rfif.rdat2[19]~256_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[24][19]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\regs[16][19]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[24][19]~q ),
	.datad(\regs[16][19]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~256_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~256 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[19]~256 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \rfif.rdat2[19]~257 (
// Equation(s):
// \rfif.rdat2[19]~257_combout  = (Instr_IF_18 & ((\rfif.rdat2[19]~256_combout  & (\regs[28][19]~q )) # (!\rfif.rdat2[19]~256_combout  & ((\regs[20][19]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[19]~256_combout ))))

	.dataa(\regs[28][19]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[20][19]~q ),
	.datad(\rfif.rdat2[19]~256_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~257_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~257 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[19]~257 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[19]~258 (
// Equation(s):
// \rfif.rdat2[19]~258_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\rfif.rdat2[19]~255_combout )))) # (!Instr_IF_16 & (!Instr_IF_17 & ((\rfif.rdat2[19]~257_combout ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[19]~255_combout ),
	.datad(\rfif.rdat2[19]~257_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~258_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~258 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[19]~258 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N20
cycloneive_lcell_comb \rfif.rdat2[19]~261 (
// Equation(s):
// \rfif.rdat2[19]~261_combout  = (Instr_IF_17 & ((\rfif.rdat2[19]~258_combout  & ((\rfif.rdat2[19]~260_combout ))) # (!\rfif.rdat2[19]~258_combout  & (\rfif.rdat2[19]~253_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[19]~258_combout ))))

	.dataa(\rfif.rdat2[19]~253_combout ),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[19]~260_combout ),
	.datad(\rfif.rdat2[19]~258_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[19]~261_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[19]~261 .lut_mask = 16'hF388;
defparam \rfif.rdat2[19]~261 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N25
dffeas \regs[21][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][18] .is_wysiwyg = "true";
defparam \regs[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N19
dffeas \regs[29][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][18] .is_wysiwyg = "true";
defparam \regs[29][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N7
dffeas \regs[17][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][18] .is_wysiwyg = "true";
defparam \regs[17][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \regs[25][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][18] .is_wysiwyg = "true";
defparam \regs[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \rfif.rdat1[18]~260 (
// Equation(s):
// \rfif.rdat1[18]~260_combout  = (Instr_IF_24 & (((\regs[25][18]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][18]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][18]~q ),
	.datac(\regs[25][18]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~260_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~260 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[18]~260 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[18]~261 (
// Equation(s):
// \rfif.rdat1[18]~261_combout  = (Instr_IF_23 & ((\rfif.rdat1[18]~260_combout  & ((\regs[29][18]~q ))) # (!\rfif.rdat1[18]~260_combout  & (\regs[21][18]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[18]~260_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[21][18]~q ),
	.datac(\regs[29][18]~q ),
	.datad(\rfif.rdat1[18]~260_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~261_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~261 .lut_mask = 16'hF588;
defparam \rfif.rdat1[18]~261 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \regs[19][18]~feeder (
// Equation(s):
// \regs[19][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b12),
	.cin(gnd),
	.combout(\regs[19][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[19][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N23
dffeas \regs[19][18] (
	.clk(!CLK),
	.d(\regs[19][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][18] .is_wysiwyg = "true";
defparam \regs[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \regs[27][18]~feeder (
// Equation(s):
// \regs[27][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b12),
	.cin(gnd),
	.combout(\regs[27][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N1
dffeas \regs[27][18] (
	.clk(!CLK),
	.d(\regs[27][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][18] .is_wysiwyg = "true";
defparam \regs[27][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[18]~267 (
// Equation(s):
// \rfif.rdat1[18]~267_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][18]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & (\regs[19][18]~q )))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[19][18]~q ),
	.datad(\regs[27][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~267_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~267 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[18]~267 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N19
dffeas \regs[23][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][18] .is_wysiwyg = "true";
defparam \regs[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N21
dffeas \regs[31][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][18] .is_wysiwyg = "true";
defparam \regs[31][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N18
cycloneive_lcell_comb \rfif.rdat1[18]~268 (
// Equation(s):
// \rfif.rdat1[18]~268_combout  = (\rfif.rdat1[18]~267_combout  & (((\regs[31][18]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[18]~267_combout  & (Instr_IF_23 & (\regs[23][18]~q )))

	.dataa(\rfif.rdat1[18]~267_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[23][18]~q ),
	.datad(\regs[31][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~268_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~268 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[18]~268 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N21
dffeas \regs[24][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][18] .is_wysiwyg = "true";
defparam \regs[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N13
dffeas \regs[20][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][18] .is_wysiwyg = "true";
defparam \regs[20][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[18]~264 (
// Equation(s):
// \rfif.rdat1[18]~264_combout  = (Instr_IF_23 & (((\regs[20][18]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][18]~q  & ((!Instr_IF_24))))

	.dataa(\regs[16][18]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][18]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~264_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~264 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[18]~264 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[18]~265 (
// Equation(s):
// \rfif.rdat1[18]~265_combout  = (Instr_IF_24 & ((\rfif.rdat1[18]~264_combout  & (\regs[28][18]~q )) # (!\rfif.rdat1[18]~264_combout  & ((\regs[24][18]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[18]~264_combout ))))

	.dataa(\regs[28][18]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[24][18]~q ),
	.datad(\rfif.rdat1[18]~264_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~265_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~265 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[18]~265 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \regs[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][18] .is_wysiwyg = "true";
defparam \regs[26][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N5
dffeas \regs[22][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][18] .is_wysiwyg = "true";
defparam \regs[22][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[18]~262 (
// Equation(s):
// \rfif.rdat1[18]~262_combout  = (Instr_IF_23 & (((\regs[22][18]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[18][18]~q  & ((!Instr_IF_24))))

	.dataa(\regs[18][18]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[22][18]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~262_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~262 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[18]~262 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[18]~263 (
// Equation(s):
// \rfif.rdat1[18]~263_combout  = (Instr_IF_24 & ((\rfif.rdat1[18]~262_combout  & (\regs[30][18]~q )) # (!\rfif.rdat1[18]~262_combout  & ((\regs[26][18]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[18]~262_combout ))))

	.dataa(\regs[30][18]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[26][18]~q ),
	.datad(\rfif.rdat1[18]~262_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~263_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~263 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[18]~263 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[18]~266 (
// Equation(s):
// \rfif.rdat1[18]~266_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[18]~263_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[18]~265_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[18]~265_combout ),
	.datad(\rfif.rdat1[18]~263_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~266_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~266 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[18]~266 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N29
dffeas \regs[15][18] (
	.clk(!CLK),
	.d(input_b12),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][18] .is_wysiwyg = "true";
defparam \regs[15][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \regs[14][18]~feeder (
// Equation(s):
// \regs[14][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b12),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][18]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N9
dffeas \regs[14][18] (
	.clk(!CLK),
	.d(\regs[14][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][18] .is_wysiwyg = "true";
defparam \regs[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \regs[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][18] .is_wysiwyg = "true";
defparam \regs[12][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \regs[13][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][18] .is_wysiwyg = "true";
defparam \regs[13][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \rfif.rdat1[18]~277 (
// Equation(s):
// \rfif.rdat1[18]~277_combout  = (Instr_IF_21 & (((\regs[13][18]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][18]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][18]~q ),
	.datac(\regs[13][18]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~277_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~277 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[18]~277 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[18]~278 (
// Equation(s):
// \rfif.rdat1[18]~278_combout  = (Instr_IF_22 & ((\rfif.rdat1[18]~277_combout  & (\regs[15][18]~q )) # (!\rfif.rdat1[18]~277_combout  & ((\regs[14][18]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[18]~277_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[15][18]~q ),
	.datac(\regs[14][18]~q ),
	.datad(\rfif.rdat1[18]~277_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~278_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~278 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[18]~278 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N19
dffeas \regs[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][18] .is_wysiwyg = "true";
defparam \regs[7][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N19
dffeas \regs[6][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][18] .is_wysiwyg = "true";
defparam \regs[6][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N21
dffeas \regs[5][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][18] .is_wysiwyg = "true";
defparam \regs[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \rfif.rdat1[18]~270 (
// Equation(s):
// \rfif.rdat1[18]~270_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][18]~q ))) # (!Instr_IF_21 & (\regs[4][18]~q ))))

	.dataa(\regs[4][18]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][18]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~270_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~270 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[18]~270 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \rfif.rdat1[18]~271 (
// Equation(s):
// \rfif.rdat1[18]~271_combout  = (Instr_IF_22 & ((\rfif.rdat1[18]~270_combout  & (\regs[7][18]~q )) # (!\rfif.rdat1[18]~270_combout  & ((\regs[6][18]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[18]~270_combout ))))

	.dataa(\regs[7][18]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[6][18]~q ),
	.datad(\rfif.rdat1[18]~270_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~271_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~271 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[18]~271 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \regs[11][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][18] .is_wysiwyg = "true";
defparam \regs[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N7
dffeas \regs[9][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][18] .is_wysiwyg = "true";
defparam \regs[9][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \regs[10][18]~feeder (
// Equation(s):
// \regs[10][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b12),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][18]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N21
dffeas \regs[10][18] (
	.clk(!CLK),
	.d(\regs[10][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][18] .is_wysiwyg = "true";
defparam \regs[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[18]~272 (
// Equation(s):
// \rfif.rdat1[18]~272_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[10][18]~q ))) # (!Instr_IF_22 & (\regs[8][18]~q ))))

	.dataa(\regs[8][18]~q ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\regs[10][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~272_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~272 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[18]~272 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \rfif.rdat1[18]~273 (
// Equation(s):
// \rfif.rdat1[18]~273_combout  = (Instr_IF_21 & ((\rfif.rdat1[18]~272_combout  & (\regs[11][18]~q )) # (!\rfif.rdat1[18]~272_combout  & ((\regs[9][18]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[18]~272_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][18]~q ),
	.datac(\regs[9][18]~q ),
	.datad(\rfif.rdat1[18]~272_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~273_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~273 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[18]~273 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \regs[1][18]~feeder (
// Equation(s):
// \regs[1][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b12),
	.cin(gnd),
	.combout(\regs[1][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N1
dffeas \regs[1][18] (
	.clk(!CLK),
	.d(\regs[1][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][18] .is_wysiwyg = "true";
defparam \regs[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \regs[3][18]~feeder (
// Equation(s):
// \regs[3][18]~feeder_combout  = \input_b~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b12),
	.cin(gnd),
	.combout(\regs[3][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][18]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N27
dffeas \regs[3][18] (
	.clk(!CLK),
	.d(\regs[3][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][18] .is_wysiwyg = "true";
defparam \regs[3][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N19
dffeas \regs[2][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][18] .is_wysiwyg = "true";
defparam \regs[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N17
dffeas \regs[0][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][18] .is_wysiwyg = "true";
defparam \regs[0][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[18]~274 (
// Equation(s):
// \rfif.rdat1[18]~274_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[2][18]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[0][18]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[2][18]~q ),
	.datad(\regs[0][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~274_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~274 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[18]~274 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[18]~275 (
// Equation(s):
// \rfif.rdat1[18]~275_combout  = (Instr_IF_21 & ((\rfif.rdat1[18]~274_combout  & ((\regs[3][18]~q ))) # (!\rfif.rdat1[18]~274_combout  & (\regs[1][18]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[18]~274_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[1][18]~q ),
	.datac(\regs[3][18]~q ),
	.datad(\rfif.rdat1[18]~274_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~275_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~275 .lut_mask = 16'hF588;
defparam \rfif.rdat1[18]~275 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[18]~276 (
// Equation(s):
// \rfif.rdat1[18]~276_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\rfif.rdat1[18]~273_combout )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\rfif.rdat1[18]~275_combout ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[18]~273_combout ),
	.datad(\rfif.rdat1[18]~275_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[18]~276_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[18]~276 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[18]~276 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[18]~274 (
// Equation(s):
// \rfif.rdat2[18]~274_combout  = (\rfif.rdat2[18]~273_combout  & (((\regs[29][18]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[18]~273_combout  & (Instr_IF_18 & (\regs[21][18]~q )))

	.dataa(\rfif.rdat2[18]~273_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[21][18]~q ),
	.datad(\regs[29][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~274_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~274 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[18]~274 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \rfif.rdat2[18]~280 (
// Equation(s):
// \rfif.rdat2[18]~280_combout  = (Instr_IF_19 & (((Instr_IF_18) # (\regs[27][18]~q )))) # (!Instr_IF_19 & (\regs[19][18]~q  & (!Instr_IF_18)))

	.dataa(\regs[19][18]~q ),
	.datab(Instr_IF_19),
	.datac(Instr_IF_18),
	.datad(\regs[27][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~280_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~280 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[18]~280 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N20
cycloneive_lcell_comb \rfif.rdat2[18]~281 (
// Equation(s):
// \rfif.rdat2[18]~281_combout  = (Instr_IF_18 & ((\rfif.rdat2[18]~280_combout  & ((\regs[31][18]~q ))) # (!\rfif.rdat2[18]~280_combout  & (\regs[23][18]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[18]~280_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][18]~q ),
	.datac(\regs[31][18]~q ),
	.datad(\rfif.rdat2[18]~280_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~281_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~281 .lut_mask = 16'hF588;
defparam \rfif.rdat2[18]~281 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N23
dffeas \regs[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][18] .is_wysiwyg = "true";
defparam \regs[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[18]~277 (
// Equation(s):
// \rfif.rdat2[18]~277_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][18]~q ))) # (!Instr_IF_18 & (\regs[16][18]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[16][18]~q ),
	.datad(\regs[20][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~277_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~277 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[18]~277 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N31
dffeas \regs[28][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][18] .is_wysiwyg = "true";
defparam \regs[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[18]~278 (
// Equation(s):
// \rfif.rdat2[18]~278_combout  = (Instr_IF_19 & ((\rfif.rdat2[18]~277_combout  & (\regs[28][18]~q )) # (!\rfif.rdat2[18]~277_combout  & ((\regs[24][18]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[18]~277_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[18]~277_combout ),
	.datac(\regs[28][18]~q ),
	.datad(\regs[24][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~278_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~278 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[18]~278 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N27
dffeas \regs[30][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][18] .is_wysiwyg = "true";
defparam \regs[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N23
dffeas \regs[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][18] .is_wysiwyg = "true";
defparam \regs[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \rfif.rdat2[18]~275 (
// Equation(s):
// \rfif.rdat2[18]~275_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[22][18]~q )) # (!Instr_IF_18 & ((\regs[18][18]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[22][18]~q ),
	.datac(\regs[18][18]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~275_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~275 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[18]~275 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \rfif.rdat2[18]~276 (
// Equation(s):
// \rfif.rdat2[18]~276_combout  = (Instr_IF_19 & ((\rfif.rdat2[18]~275_combout  & ((\regs[30][18]~q ))) # (!\rfif.rdat2[18]~275_combout  & (\regs[26][18]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[18]~275_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][18]~q ),
	.datac(\regs[30][18]~q ),
	.datad(\rfif.rdat2[18]~275_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~276_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~276 .lut_mask = 16'hF588;
defparam \rfif.rdat2[18]~276 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \rfif.rdat2[18]~279 (
// Equation(s):
// \rfif.rdat2[18]~279_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[18]~276_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[18]~278_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[18]~278_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[18]~276_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~279_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~279 .lut_mask = 16'hF4A4;
defparam \rfif.rdat2[18]~279 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[18]~282 (
// Equation(s):
// \rfif.rdat2[18]~282_combout  = (Instr_IF_16 & ((\rfif.rdat2[18]~279_combout  & ((\rfif.rdat2[18]~281_combout ))) # (!\rfif.rdat2[18]~279_combout  & (\rfif.rdat2[18]~274_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[18]~279_combout ))))

	.dataa(\rfif.rdat2[18]~274_combout ),
	.datab(\rfif.rdat2[18]~281_combout ),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[18]~279_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~282_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~282 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[18]~282 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N31
dffeas \regs[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][18] .is_wysiwyg = "true";
defparam \regs[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[18]~285 (
// Equation(s):
// \rfif.rdat2[18]~285_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][18]~q ))) # (!Instr_IF_17 & (\regs[8][18]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][18]~q ),
	.datad(\regs[10][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~285_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~285 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[18]~285 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[18]~286 (
// Equation(s):
// \rfif.rdat2[18]~286_combout  = (Instr_IF_16 & ((\rfif.rdat2[18]~285_combout  & (\regs[11][18]~q )) # (!\rfif.rdat2[18]~285_combout  & ((\regs[9][18]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[18]~285_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[18]~285_combout ),
	.datac(\regs[11][18]~q ),
	.datad(\regs[9][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~286_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~286 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[18]~286 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[18]~287 (
// Equation(s):
// \rfif.rdat2[18]~287_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][18]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][18]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][18]~q ),
	.datad(\regs[2][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~287_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~287 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[18]~287 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[18]~288 (
// Equation(s):
// \rfif.rdat2[18]~288_combout  = (Instr_IF_16 & ((\rfif.rdat2[18]~287_combout  & ((\regs[3][18]~q ))) # (!\rfif.rdat2[18]~287_combout  & (\regs[1][18]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[18]~287_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][18]~q ),
	.datac(\regs[3][18]~q ),
	.datad(\rfif.rdat2[18]~287_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~288_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~288 .lut_mask = 16'hF588;
defparam \rfif.rdat2[18]~288 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[18]~289 (
// Equation(s):
// \rfif.rdat2[18]~289_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[18]~286_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[18]~288_combout )))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[18]~286_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[18]~288_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~289_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~289 .lut_mask = 16'hE5E0;
defparam \rfif.rdat2[18]~289 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N9
dffeas \regs[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][18] .is_wysiwyg = "true";
defparam \regs[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \rfif.rdat2[18]~283 (
// Equation(s):
// \rfif.rdat2[18]~283_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][18]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][18]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][18]~q ),
	.datad(\regs[5][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~283_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~283 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[18]~283 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[18]~284 (
// Equation(s):
// \rfif.rdat2[18]~284_combout  = (Instr_IF_17 & ((\rfif.rdat2[18]~283_combout  & ((\regs[7][18]~q ))) # (!\rfif.rdat2[18]~283_combout  & (\regs[6][18]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[18]~283_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[6][18]~q ),
	.datac(\regs[7][18]~q ),
	.datad(\rfif.rdat2[18]~283_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~284_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~284 .lut_mask = 16'hF588;
defparam \rfif.rdat2[18]~284 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \rfif.rdat2[18]~290 (
// Equation(s):
// \rfif.rdat2[18]~290_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][18]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][18]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][18]~q ),
	.datad(\regs[13][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~290_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~290 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[18]~290 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[18]~291 (
// Equation(s):
// \rfif.rdat2[18]~291_combout  = (Instr_IF_17 & ((\rfif.rdat2[18]~290_combout  & ((\regs[15][18]~q ))) # (!\rfif.rdat2[18]~290_combout  & (\regs[14][18]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[18]~290_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[14][18]~q ),
	.datac(\rfif.rdat2[18]~290_combout ),
	.datad(\regs[15][18]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~291_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~291 .lut_mask = 16'hF858;
defparam \rfif.rdat2[18]~291 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[18]~292 (
// Equation(s):
// \rfif.rdat2[18]~292_combout  = (Instr_IF_18 & ((\rfif.rdat2[18]~289_combout  & ((\rfif.rdat2[18]~291_combout ))) # (!\rfif.rdat2[18]~289_combout  & (\rfif.rdat2[18]~284_combout )))) # (!Instr_IF_18 & (\rfif.rdat2[18]~289_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[18]~289_combout ),
	.datac(\rfif.rdat2[18]~284_combout ),
	.datad(\rfif.rdat2[18]~291_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[18]~292_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[18]~292 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[18]~292 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N19
dffeas \regs[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][17] .is_wysiwyg = "true";
defparam \regs[18][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N31
dffeas \regs[26][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][17] .is_wysiwyg = "true";
defparam \regs[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \rfif.rdat1[17]~280 (
// Equation(s):
// \rfif.rdat1[17]~280_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[26][17]~q ))) # (!Instr_IF_24 & (\regs[18][17]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[18][17]~q ),
	.datac(\regs[26][17]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~280_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~280 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[17]~280 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N5
dffeas \regs[30][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][17] .is_wysiwyg = "true";
defparam \regs[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N5
dffeas \regs[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][17] .is_wysiwyg = "true";
defparam \regs[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[17]~281 (
// Equation(s):
// \rfif.rdat1[17]~281_combout  = (\rfif.rdat1[17]~280_combout  & (((\regs[30][17]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[17]~280_combout  & (Instr_IF_23 & ((\regs[22][17]~q ))))

	.dataa(\rfif.rdat1[17]~280_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[30][17]~q ),
	.datad(\regs[22][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~281_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~281 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[17]~281 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N29
dffeas \regs[21][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][17] .is_wysiwyg = "true";
defparam \regs[21][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[17]~282 (
// Equation(s):
// \rfif.rdat1[17]~282_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][17]~q ))) # (!Instr_IF_23 & (\regs[17][17]~q ))))

	.dataa(\regs[17][17]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[21][17]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~282_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~282 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[17]~282 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas \regs[25][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][17] .is_wysiwyg = "true";
defparam \regs[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N7
dffeas \regs[29][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][17] .is_wysiwyg = "true";
defparam \regs[29][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[17]~283 (
// Equation(s):
// \rfif.rdat1[17]~283_combout  = (Instr_IF_24 & ((\rfif.rdat1[17]~282_combout  & ((\regs[29][17]~q ))) # (!\rfif.rdat1[17]~282_combout  & (\regs[25][17]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[17]~282_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[17]~282_combout ),
	.datac(\regs[25][17]~q ),
	.datad(\regs[29][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~283_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~283 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[17]~283 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N17
dffeas \regs[20][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][17] .is_wysiwyg = "true";
defparam \regs[20][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N17
dffeas \regs[28][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][17] .is_wysiwyg = "true";
defparam \regs[28][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \rfif.rdat1[17]~285 (
// Equation(s):
// \rfif.rdat1[17]~285_combout  = (\rfif.rdat1[17]~284_combout  & (((\regs[28][17]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[17]~284_combout  & (Instr_IF_23 & (\regs[20][17]~q )))

	.dataa(\rfif.rdat1[17]~284_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[20][17]~q ),
	.datad(\regs[28][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~285_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~285 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[17]~285 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \rfif.rdat1[17]~286 (
// Equation(s):
// \rfif.rdat1[17]~286_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\rfif.rdat1[17]~283_combout )) # (!Instr_IF_21 & ((\rfif.rdat1[17]~285_combout )))))

	.dataa(\rfif.rdat1[17]~283_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[17]~285_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~286_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~286 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[17]~286 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \regs[27][17]~feeder (
// Equation(s):
// \regs[27][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b13),
	.cin(gnd),
	.combout(\regs[27][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \regs[27][17] (
	.clk(!CLK),
	.d(\regs[27][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][17] .is_wysiwyg = "true";
defparam \regs[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N11
dffeas \regs[23][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][17] .is_wysiwyg = "true";
defparam \regs[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N3
dffeas \regs[19][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][17] .is_wysiwyg = "true";
defparam \regs[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N10
cycloneive_lcell_comb \rfif.rdat1[17]~287 (
// Equation(s):
// \rfif.rdat1[17]~287_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][17]~q )) # (!Instr_IF_23 & ((\regs[19][17]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][17]~q ),
	.datad(\regs[19][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~287_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~287 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[17]~287 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \regs[31][17]~feeder (
// Equation(s):
// \regs[31][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b13),
	.cin(gnd),
	.combout(\regs[31][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N3
dffeas \regs[31][17] (
	.clk(!CLK),
	.d(\regs[31][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][17] .is_wysiwyg = "true";
defparam \regs[31][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[17]~288 (
// Equation(s):
// \rfif.rdat1[17]~288_combout  = (Instr_IF_24 & ((\rfif.rdat1[17]~287_combout  & ((\regs[31][17]~q ))) # (!\rfif.rdat1[17]~287_combout  & (\regs[27][17]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[17]~287_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[27][17]~q ),
	.datac(\rfif.rdat1[17]~287_combout ),
	.datad(\regs[31][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~288_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~288 .lut_mask = 16'hF858;
defparam \rfif.rdat1[17]~288 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N13
dffeas \regs[13][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][17] .is_wysiwyg = "true";
defparam \regs[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \regs[15][17]~feeder (
// Equation(s):
// \regs[15][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b13),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][17]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N1
dffeas \regs[15][17] (
	.clk(!CLK),
	.d(\regs[15][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][17] .is_wysiwyg = "true";
defparam \regs[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N19
dffeas \regs[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][17] .is_wysiwyg = "true";
defparam \regs[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[17]~297 (
// Equation(s):
// \rfif.rdat1[17]~297_combout  = (Instr_IF_22 & ((\regs[14][17]~q ) # ((Instr_IF_21)))) # (!Instr_IF_22 & (((\regs[12][17]~q  & !Instr_IF_21))))

	.dataa(\regs[14][17]~q ),
	.datab(\regs[12][17]~q ),
	.datac(Instr_IF_22),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~297_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~297 .lut_mask = 16'hF0AC;
defparam \rfif.rdat1[17]~297 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[17]~298 (
// Equation(s):
// \rfif.rdat1[17]~298_combout  = (Instr_IF_21 & ((\rfif.rdat1[17]~297_combout  & ((\regs[15][17]~q ))) # (!\rfif.rdat1[17]~297_combout  & (\regs[13][17]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[17]~297_combout ))))

	.dataa(\regs[13][17]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[15][17]~q ),
	.datad(\rfif.rdat1[17]~297_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~298_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~298 .lut_mask = 16'hF388;
defparam \rfif.rdat1[17]~298 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N15
dffeas \regs[9][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][17] .is_wysiwyg = "true";
defparam \regs[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N9
dffeas \regs[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][17] .is_wysiwyg = "true";
defparam \regs[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[17]~290 (
// Equation(s):
// \rfif.rdat1[17]~290_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][17]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[8][17]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[9][17]~q ),
	.datad(\regs[8][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~290_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~290 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[17]~290 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N17
dffeas \regs[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][17] .is_wysiwyg = "true";
defparam \regs[11][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N15
dffeas \regs[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][17] .is_wysiwyg = "true";
defparam \regs[10][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[17]~291 (
// Equation(s):
// \rfif.rdat1[17]~291_combout  = (Instr_IF_22 & ((\rfif.rdat1[17]~290_combout  & (\regs[11][17]~q )) # (!\rfif.rdat1[17]~290_combout  & ((\regs[10][17]~q ))))) # (!Instr_IF_22 & (\rfif.rdat1[17]~290_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[17]~290_combout ),
	.datac(\regs[11][17]~q ),
	.datad(\regs[10][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~291_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~291 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[17]~291 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N5
dffeas \regs[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][17] .is_wysiwyg = "true";
defparam \regs[1][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N1
dffeas \regs[0][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][17] .is_wysiwyg = "true";
defparam \regs[0][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[17]~294 (
// Equation(s):
// \rfif.rdat1[17]~294_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][17]~q )) # (!Instr_IF_21 & ((\regs[0][17]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][17]~q ),
	.datad(\regs[0][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~294_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~294 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[17]~294 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \regs[3][17]~feeder (
// Equation(s):
// \regs[3][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b13),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][17]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N9
dffeas \regs[3][17] (
	.clk(!CLK),
	.d(\regs[3][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][17] .is_wysiwyg = "true";
defparam \regs[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[17]~295 (
// Equation(s):
// \rfif.rdat1[17]~295_combout  = (\rfif.rdat1[17]~294_combout  & (((\regs[3][17]~q ) # (!Instr_IF_22)))) # (!\rfif.rdat1[17]~294_combout  & (\regs[2][17]~q  & (Instr_IF_22)))

	.dataa(\regs[2][17]~q ),
	.datab(\rfif.rdat1[17]~294_combout ),
	.datac(Instr_IF_22),
	.datad(\regs[3][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~295_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~295 .lut_mask = 16'hEC2C;
defparam \rfif.rdat1[17]~295 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N3
dffeas \regs[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][17] .is_wysiwyg = "true";
defparam \regs[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N25
dffeas \regs[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][17] .is_wysiwyg = "true";
defparam \regs[5][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[17]~293 (
// Equation(s):
// \rfif.rdat1[17]~293_combout  = (\rfif.rdat1[17]~292_combout  & ((\regs[7][17]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[17]~292_combout  & (((\regs[5][17]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[17]~292_combout ),
	.datab(\regs[7][17]~q ),
	.datac(\regs[5][17]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~293_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~293 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[17]~293 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[17]~296 (
// Equation(s):
// \rfif.rdat1[17]~296_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\rfif.rdat1[17]~293_combout )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\rfif.rdat1[17]~295_combout )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[17]~295_combout ),
	.datad(\rfif.rdat1[17]~293_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[17]~296_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[17]~296 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[17]~296 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N23
dffeas \regs[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][17] .is_wysiwyg = "true";
defparam \regs[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[17]~296 (
// Equation(s):
// \rfif.rdat2[17]~296_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][17]~q ))) # (!Instr_IF_18 & (\regs[17][17]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][17]~q ),
	.datad(\regs[21][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~296_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~296 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[17]~296 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[17]~297 (
// Equation(s):
// \rfif.rdat2[17]~297_combout  = (\rfif.rdat2[17]~296_combout  & (((\regs[29][17]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[17]~296_combout  & (\regs[25][17]~q  & ((Instr_IF_19))))

	.dataa(\regs[25][17]~q ),
	.datab(\rfif.rdat2[17]~296_combout ),
	.datac(\regs[29][17]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~297_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~297 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[17]~297 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N2
cycloneive_lcell_comb \regs[24][17]~feeder (
// Equation(s):
// \regs[24][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b13),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[24][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[24][17]~feeder .lut_mask = 16'hF0F0;
defparam \regs[24][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N3
dffeas \regs[24][17] (
	.clk(!CLK),
	.d(\regs[24][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][17] .is_wysiwyg = "true";
defparam \regs[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[17]~298 (
// Equation(s):
// \rfif.rdat2[17]~298_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][17]~q ))) # (!Instr_IF_19 & (\regs[16][17]~q ))))

	.dataa(\regs[16][17]~q ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\regs[24][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~298_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~298 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[17]~298 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[17]~299 (
// Equation(s):
// \rfif.rdat2[17]~299_combout  = (Instr_IF_18 & ((\rfif.rdat2[17]~298_combout  & ((\regs[28][17]~q ))) # (!\rfif.rdat2[17]~298_combout  & (\regs[20][17]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[17]~298_combout ))))

	.dataa(\regs[20][17]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][17]~q ),
	.datad(\rfif.rdat2[17]~298_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~299_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~299 .lut_mask = 16'hF388;
defparam \rfif.rdat2[17]~299 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[17]~300 (
// Equation(s):
// \rfif.rdat2[17]~300_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[17]~297_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[17]~299_combout )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[17]~297_combout ),
	.datad(\rfif.rdat2[17]~299_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~300_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~300 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[17]~300 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[17]~301 (
// Equation(s):
// \rfif.rdat2[17]~301_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[23][17]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[19][17]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][17]~q ),
	.datad(\regs[23][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~301_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~301 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[17]~301 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[17]~302 (
// Equation(s):
// \rfif.rdat2[17]~302_combout  = (Instr_IF_19 & ((\rfif.rdat2[17]~301_combout  & (\regs[31][17]~q )) # (!\rfif.rdat2[17]~301_combout  & ((\regs[27][17]~q ))))) # (!Instr_IF_19 & (((\rfif.rdat2[17]~301_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[31][17]~q ),
	.datac(\rfif.rdat2[17]~301_combout ),
	.datad(\regs[27][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~302_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~302 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[17]~302 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[17]~294 (
// Equation(s):
// \rfif.rdat2[17]~294_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][17]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][17]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][17]~q ),
	.datad(\regs[26][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~294_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~294 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[17]~294 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[17]~295 (
// Equation(s):
// \rfif.rdat2[17]~295_combout  = (Instr_IF_18 & ((\rfif.rdat2[17]~294_combout  & (\regs[30][17]~q )) # (!\rfif.rdat2[17]~294_combout  & ((\regs[22][17]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[17]~294_combout ))))

	.dataa(\regs[30][17]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][17]~q ),
	.datad(\rfif.rdat2[17]~294_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~295_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~295 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[17]~295 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[17]~303 (
// Equation(s):
// \rfif.rdat2[17]~303_combout  = (\rfif.rdat2[17]~300_combout  & ((\rfif.rdat2[17]~302_combout ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[17]~300_combout  & (((\rfif.rdat2[17]~295_combout  & Instr_IF_17))))

	.dataa(\rfif.rdat2[17]~300_combout ),
	.datab(\rfif.rdat2[17]~302_combout ),
	.datac(\rfif.rdat2[17]~295_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~303_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~303 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[17]~303 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \rfif.rdat2[17]~304 (
// Equation(s):
// \rfif.rdat2[17]~304_combout  = (Instr_IF_16 & ((\regs[9][17]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[8][17]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][17]~q ),
	.datac(\regs[8][17]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~304_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~304 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[17]~304 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \rfif.rdat2[17]~305 (
// Equation(s):
// \rfif.rdat2[17]~305_combout  = (Instr_IF_17 & ((\rfif.rdat2[17]~304_combout  & ((\regs[11][17]~q ))) # (!\rfif.rdat2[17]~304_combout  & (\regs[10][17]~q )))) # (!Instr_IF_17 & (\rfif.rdat2[17]~304_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[17]~304_combout ),
	.datac(\regs[10][17]~q ),
	.datad(\regs[11][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~305_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~305 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[17]~305 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \regs[14][17]~feeder (
// Equation(s):
// \regs[14][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b13),
	.cin(gnd),
	.combout(\regs[14][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][17]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N23
dffeas \regs[14][17] (
	.clk(!CLK),
	.d(\regs[14][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][17] .is_wysiwyg = "true";
defparam \regs[14][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \rfif.rdat2[17]~311 (
// Equation(s):
// \rfif.rdat2[17]~311_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[14][17]~q )) # (!Instr_IF_17 & ((\regs[12][17]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[14][17]~q ),
	.datac(\regs[12][17]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~311_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~311 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[17]~311 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \rfif.rdat2[17]~312 (
// Equation(s):
// \rfif.rdat2[17]~312_combout  = (Instr_IF_16 & ((\rfif.rdat2[17]~311_combout  & ((\regs[15][17]~q ))) # (!\rfif.rdat2[17]~311_combout  & (\regs[13][17]~q )))) # (!Instr_IF_16 & (\rfif.rdat2[17]~311_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[17]~311_combout ),
	.datac(\regs[13][17]~q ),
	.datad(\regs[15][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~312_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~312 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[17]~312 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N19
dffeas \regs[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][17] .is_wysiwyg = "true";
defparam \regs[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \regs[6][17]~feeder (
// Equation(s):
// \regs[6][17]~feeder_combout  = \input_b~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b13),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[6][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][17]~feeder .lut_mask = 16'hF0F0;
defparam \regs[6][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N29
dffeas \regs[6][17] (
	.clk(!CLK),
	.d(\regs[6][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][17] .is_wysiwyg = "true";
defparam \regs[6][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[17]~306 (
// Equation(s):
// \rfif.rdat2[17]~306_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][17]~q ))) # (!Instr_IF_17 & (\regs[4][17]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][17]~q ),
	.datad(\regs[6][17]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~306_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~306 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[17]~306 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[17]~307 (
// Equation(s):
// \rfif.rdat2[17]~307_combout  = (Instr_IF_16 & ((\rfif.rdat2[17]~306_combout  & ((\regs[7][17]~q ))) # (!\rfif.rdat2[17]~306_combout  & (\regs[5][17]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[17]~306_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][17]~q ),
	.datac(\regs[7][17]~q ),
	.datad(\rfif.rdat2[17]~306_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~307_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~307 .lut_mask = 16'hF588;
defparam \rfif.rdat2[17]~307 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \rfif.rdat2[17]~310 (
// Equation(s):
// \rfif.rdat2[17]~310_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & ((\rfif.rdat2[17]~307_combout ))) # (!Instr_IF_18 & (\rfif.rdat2[17]~309_combout ))))

	.dataa(\rfif.rdat2[17]~309_combout ),
	.datab(Instr_IF_19),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[17]~307_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~310_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~310 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[17]~310 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[17]~313 (
// Equation(s):
// \rfif.rdat2[17]~313_combout  = (\rfif.rdat2[17]~310_combout  & (((\rfif.rdat2[17]~312_combout ) # (!Instr_IF_19)))) # (!\rfif.rdat2[17]~310_combout  & (\rfif.rdat2[17]~305_combout  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[17]~305_combout ),
	.datab(\rfif.rdat2[17]~312_combout ),
	.datac(\rfif.rdat2[17]~310_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[17]~313_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[17]~313 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[17]~313 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N3
dffeas \regs[31][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][16] .is_wysiwyg = "true";
defparam \regs[31][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N29
dffeas \regs[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][16] .is_wysiwyg = "true";
defparam \regs[23][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N26
cycloneive_lcell_comb \regs[27][16]~feeder (
// Equation(s):
// \regs[27][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b14),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N27
dffeas \regs[27][16] (
	.clk(!CLK),
	.d(\regs[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][16] .is_wysiwyg = "true";
defparam \regs[27][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \regs[19][16]~feeder (
// Equation(s):
// \regs[19][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b14),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[19][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[19][16]~feeder .lut_mask = 16'hF0F0;
defparam \regs[19][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N25
dffeas \regs[19][16] (
	.clk(!CLK),
	.d(\regs[19][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][16] .is_wysiwyg = "true";
defparam \regs[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N12
cycloneive_lcell_comb \rfif.rdat1[16]~307 (
// Equation(s):
// \rfif.rdat1[16]~307_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[27][16]~q )) # (!Instr_IF_24 & ((\regs[19][16]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[27][16]~q ),
	.datad(\regs[19][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~307_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~307 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[16]~307 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N28
cycloneive_lcell_comb \rfif.rdat1[16]~308 (
// Equation(s):
// \rfif.rdat1[16]~308_combout  = (Instr_IF_23 & ((\rfif.rdat1[16]~307_combout  & (\regs[31][16]~q )) # (!\rfif.rdat1[16]~307_combout  & ((\regs[23][16]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[16]~307_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[31][16]~q ),
	.datac(\regs[23][16]~q ),
	.datad(\rfif.rdat1[16]~307_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~308_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~308 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[16]~308 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N1
dffeas \regs[24][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][16] .is_wysiwyg = "true";
defparam \regs[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N23
dffeas \regs[28][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][16] .is_wysiwyg = "true";
defparam \regs[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[16]~305 (
// Equation(s):
// \rfif.rdat1[16]~305_combout  = (\rfif.rdat1[16]~304_combout  & (((\regs[28][16]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[16]~304_combout  & (Instr_IF_24 & (\regs[24][16]~q )))

	.dataa(\rfif.rdat1[16]~304_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[24][16]~q ),
	.datad(\regs[28][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~305_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~305 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[16]~305 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N17
dffeas \regs[26][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][16] .is_wysiwyg = "true";
defparam \regs[26][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N19
dffeas \regs[30][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][16] .is_wysiwyg = "true";
defparam \regs[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \rfif.rdat1[16]~303 (
// Equation(s):
// \rfif.rdat1[16]~303_combout  = (\rfif.rdat1[16]~302_combout  & (((\regs[30][16]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[16]~302_combout  & (Instr_IF_24 & (\regs[26][16]~q )))

	.dataa(\rfif.rdat1[16]~302_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[26][16]~q ),
	.datad(\regs[30][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~303_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~303 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[16]~303 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \rfif.rdat1[16]~306 (
// Equation(s):
// \rfif.rdat1[16]~306_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[16]~303_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[16]~305_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[16]~305_combout ),
	.datad(\rfif.rdat1[16]~303_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~306_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~306 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[16]~306 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N5
dffeas \regs[25][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][16] .is_wysiwyg = "true";
defparam \regs[25][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N15
dffeas \regs[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][16] .is_wysiwyg = "true";
defparam \regs[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[16]~300 (
// Equation(s):
// \rfif.rdat1[16]~300_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[25][16]~q )) # (!Instr_IF_24 & ((\regs[17][16]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[25][16]~q ),
	.datad(\regs[17][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~300_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~300 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[16]~300 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \regs[29][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][16] .is_wysiwyg = "true";
defparam \regs[29][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N5
dffeas \regs[21][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][16] .is_wysiwyg = "true";
defparam \regs[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[16]~301 (
// Equation(s):
// \rfif.rdat1[16]~301_combout  = (Instr_IF_23 & ((\rfif.rdat1[16]~300_combout  & (\regs[29][16]~q )) # (!\rfif.rdat1[16]~300_combout  & ((\regs[21][16]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[16]~300_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[16]~300_combout ),
	.datac(\regs[29][16]~q ),
	.datad(\regs[21][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~301_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~301 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[16]~301 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N7
dffeas \regs[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][16] .is_wysiwyg = "true";
defparam \regs[10][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N17
dffeas \regs[8][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][16] .is_wysiwyg = "true";
defparam \regs[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \rfif.rdat1[16]~312 (
// Equation(s):
// \rfif.rdat1[16]~312_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[10][16]~q )) # (!Instr_IF_22 & ((\regs[8][16]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[10][16]~q ),
	.datad(\regs[8][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~312_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~312 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[16]~312 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N1
dffeas \regs[9][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][16] .is_wysiwyg = "true";
defparam \regs[9][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \rfif.rdat1[16]~313 (
// Equation(s):
// \rfif.rdat1[16]~313_combout  = (\rfif.rdat1[16]~312_combout  & ((\regs[11][16]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[16]~312_combout  & (((\regs[9][16]~q  & Instr_IF_21))))

	.dataa(\regs[11][16]~q ),
	.datab(\rfif.rdat1[16]~312_combout ),
	.datac(\regs[9][16]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~313_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~313 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[16]~313 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \regs[1][16]~feeder (
// Equation(s):
// \regs[1][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b14),
	.cin(gnd),
	.combout(\regs[1][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N29
dffeas \regs[1][16] (
	.clk(!CLK),
	.d(\regs[1][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][16] .is_wysiwyg = "true";
defparam \regs[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \regs[2][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][16] .is_wysiwyg = "true";
defparam \regs[2][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[16]~314 (
// Equation(s):
// \rfif.rdat1[16]~314_combout  = (Instr_IF_22 & (((\regs[2][16]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[0][16]~q  & ((!Instr_IF_21))))

	.dataa(\regs[0][16]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[2][16]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~314_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~314 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[16]~314 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[16]~315 (
// Equation(s):
// \rfif.rdat1[16]~315_combout  = (Instr_IF_21 & ((\rfif.rdat1[16]~314_combout  & (\regs[3][16]~q )) # (!\rfif.rdat1[16]~314_combout  & ((\regs[1][16]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[16]~314_combout ))))

	.dataa(\regs[3][16]~q ),
	.datab(\regs[1][16]~q ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[16]~314_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~315_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~315 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[16]~315 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \rfif.rdat1[16]~316 (
// Equation(s):
// \rfif.rdat1[16]~316_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\rfif.rdat1[16]~313_combout )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\rfif.rdat1[16]~315_combout ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[16]~313_combout ),
	.datad(\rfif.rdat1[16]~315_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~316_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~316 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[16]~316 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N7
dffeas \regs[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][16] .is_wysiwyg = "true";
defparam \regs[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N27
dffeas \regs[6][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][16] .is_wysiwyg = "true";
defparam \regs[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N17
dffeas \regs[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][16] .is_wysiwyg = "true";
defparam \regs[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[16]~310 (
// Equation(s):
// \rfif.rdat1[16]~310_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][16]~q ))) # (!Instr_IF_21 & (\regs[4][16]~q ))))

	.dataa(\regs[4][16]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][16]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~310_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~310 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[16]~310 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \rfif.rdat1[16]~311 (
// Equation(s):
// \rfif.rdat1[16]~311_combout  = (Instr_IF_22 & ((\rfif.rdat1[16]~310_combout  & (\regs[7][16]~q )) # (!\rfif.rdat1[16]~310_combout  & ((\regs[6][16]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[16]~310_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[7][16]~q ),
	.datac(\regs[6][16]~q ),
	.datad(\rfif.rdat1[16]~310_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~311_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~311 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[16]~311 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \regs[15][16]~feeder (
// Equation(s):
// \regs[15][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b14),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][16]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N7
dffeas \regs[15][16] (
	.clk(!CLK),
	.d(\regs[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][16] .is_wysiwyg = "true";
defparam \regs[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \regs[13][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][16] .is_wysiwyg = "true";
defparam \regs[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \rfif.rdat1[16]~317 (
// Equation(s):
// \rfif.rdat1[16]~317_combout  = (Instr_IF_21 & (((\regs[13][16]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][16]~q  & ((!Instr_IF_22))))

	.dataa(\regs[12][16]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][16]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~317_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~317 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[16]~317 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \regs[14][16]~feeder (
// Equation(s):
// \regs[14][16]~feeder_combout  = \input_b~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b14),
	.cin(gnd),
	.combout(\regs[14][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][16]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N15
dffeas \regs[14][16] (
	.clk(!CLK),
	.d(\regs[14][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][16] .is_wysiwyg = "true";
defparam \regs[14][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[16]~318 (
// Equation(s):
// \rfif.rdat1[16]~318_combout  = (Instr_IF_22 & ((\rfif.rdat1[16]~317_combout  & (\regs[15][16]~q )) # (!\rfif.rdat1[16]~317_combout  & ((\regs[14][16]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[16]~317_combout ))))

	.dataa(\regs[15][16]~q ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[16]~317_combout ),
	.datad(\regs[14][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[16]~318_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[16]~318 .lut_mask = 16'hBCB0;
defparam \rfif.rdat1[16]~318 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N31
dffeas \regs[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][16] .is_wysiwyg = "true";
defparam \regs[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \rfif.rdat2[16]~332 (
// Equation(s):
// \rfif.rdat2[16]~332_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][16]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][16]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][16]~q ),
	.datad(\regs[13][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~332_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~332 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[16]~332 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[16]~333 (
// Equation(s):
// \rfif.rdat2[16]~333_combout  = (Instr_IF_17 & ((\rfif.rdat2[16]~332_combout  & (\regs[15][16]~q )) # (!\rfif.rdat2[16]~332_combout  & ((\regs[14][16]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[16]~332_combout ))))

	.dataa(\regs[15][16]~q ),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[16]~332_combout ),
	.datad(\regs[14][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~333_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~333 .lut_mask = 16'hBCB0;
defparam \rfif.rdat2[16]~333 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N27
dffeas \regs[0][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][16] .is_wysiwyg = "true";
defparam \regs[0][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[16]~329 (
// Equation(s):
// \rfif.rdat2[16]~329_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][16]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][16]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][16]~q ),
	.datad(\regs[2][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~329_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~329 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[16]~329 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[16]~330 (
// Equation(s):
// \rfif.rdat2[16]~330_combout  = (Instr_IF_16 & ((\rfif.rdat2[16]~329_combout  & (\regs[3][16]~q )) # (!\rfif.rdat2[16]~329_combout  & ((\regs[1][16]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[16]~329_combout ))))

	.dataa(\regs[3][16]~q ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[16]~329_combout ),
	.datad(\regs[1][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~330_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~330 .lut_mask = 16'hBCB0;
defparam \rfif.rdat2[16]~330 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N27
dffeas \regs[11][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][16] .is_wysiwyg = "true";
defparam \regs[11][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[16]~328 (
// Equation(s):
// \rfif.rdat2[16]~328_combout  = (\rfif.rdat2[16]~327_combout  & (((\regs[11][16]~q )) # (!Instr_IF_16))) # (!\rfif.rdat2[16]~327_combout  & (Instr_IF_16 & ((\regs[9][16]~q ))))

	.dataa(\rfif.rdat2[16]~327_combout ),
	.datab(Instr_IF_16),
	.datac(\regs[11][16]~q ),
	.datad(\regs[9][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~328_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~328 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[16]~328 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[16]~331 (
// Equation(s):
// \rfif.rdat2[16]~331_combout  = (Instr_IF_19 & (((Instr_IF_18) # (\rfif.rdat2[16]~328_combout )))) # (!Instr_IF_19 & (\rfif.rdat2[16]~330_combout  & (!Instr_IF_18)))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[16]~330_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[16]~328_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~331_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~331 .lut_mask = 16'hAEA4;
defparam \rfif.rdat2[16]~331 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N9
dffeas \regs[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][16] .is_wysiwyg = "true";
defparam \regs[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \rfif.rdat2[16]~325 (
// Equation(s):
// \rfif.rdat2[16]~325_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[5][16]~q )) # (!Instr_IF_16 & ((\regs[4][16]~q )))))

	.dataa(\regs[5][16]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[4][16]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~325_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~325 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[16]~325 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[16]~326 (
// Equation(s):
// \rfif.rdat2[16]~326_combout  = (Instr_IF_17 & ((\rfif.rdat2[16]~325_combout  & (\regs[7][16]~q )) # (!\rfif.rdat2[16]~325_combout  & ((\regs[6][16]~q ))))) # (!Instr_IF_17 & (\rfif.rdat2[16]~325_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[16]~325_combout ),
	.datac(\regs[7][16]~q ),
	.datad(\regs[6][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~326_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~326 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[16]~326 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[16]~334 (
// Equation(s):
// \rfif.rdat2[16]~334_combout  = (Instr_IF_18 & ((\rfif.rdat2[16]~331_combout  & (\rfif.rdat2[16]~333_combout )) # (!\rfif.rdat2[16]~331_combout  & ((\rfif.rdat2[16]~326_combout ))))) # (!Instr_IF_18 & (((\rfif.rdat2[16]~331_combout ))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[16]~333_combout ),
	.datac(\rfif.rdat2[16]~331_combout ),
	.datad(\rfif.rdat2[16]~326_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~334_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~334 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[16]~334 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \rfif.rdat2[16]~322 (
// Equation(s):
// \rfif.rdat2[16]~322_combout  = (Instr_IF_19 & ((\regs[27][16]~q ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((!Instr_IF_18 & \regs[19][16]~q ))))

	.dataa(\regs[27][16]~q ),
	.datab(Instr_IF_19),
	.datac(Instr_IF_18),
	.datad(\regs[19][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~322_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~322 .lut_mask = 16'hCBC8;
defparam \rfif.rdat2[16]~322 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N2
cycloneive_lcell_comb \rfif.rdat2[16]~323 (
// Equation(s):
// \rfif.rdat2[16]~323_combout  = (Instr_IF_18 & ((\rfif.rdat2[16]~322_combout  & ((\regs[31][16]~q ))) # (!\rfif.rdat2[16]~322_combout  & (\regs[23][16]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[16]~322_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][16]~q ),
	.datac(\regs[31][16]~q ),
	.datad(\rfif.rdat2[16]~322_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~323_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~323 .lut_mask = 16'hF588;
defparam \rfif.rdat2[16]~323 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[16]~320 (
// Equation(s):
// \rfif.rdat2[16]~320_combout  = (\rfif.rdat2[16]~319_combout  & (((\regs[28][16]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[16]~319_combout  & (\regs[24][16]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[16]~319_combout ),
	.datab(\regs[24][16]~q ),
	.datac(\regs[28][16]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~320_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~320 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[16]~320 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \rfif.rdat2[16]~321 (
// Equation(s):
// \rfif.rdat2[16]~321_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\rfif.rdat2[16]~318_combout )) # (!Instr_IF_17 & ((\rfif.rdat2[16]~320_combout )))))

	.dataa(\rfif.rdat2[16]~318_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[16]~320_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~321_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~321 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[16]~321 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[16]~315 (
// Equation(s):
// \rfif.rdat2[16]~315_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[25][16]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[17][16]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][16]~q ),
	.datad(\regs[25][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~315_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~315 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[16]~315 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \rfif.rdat2[16]~316 (
// Equation(s):
// \rfif.rdat2[16]~316_combout  = (Instr_IF_18 & ((\rfif.rdat2[16]~315_combout  & ((\regs[29][16]~q ))) # (!\rfif.rdat2[16]~315_combout  & (\regs[21][16]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[16]~315_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[16]~315_combout ),
	.datac(\regs[21][16]~q ),
	.datad(\regs[29][16]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~316_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~316 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[16]~316 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[16]~324 (
// Equation(s):
// \rfif.rdat2[16]~324_combout  = (Instr_IF_16 & ((\rfif.rdat2[16]~321_combout  & (\rfif.rdat2[16]~323_combout )) # (!\rfif.rdat2[16]~321_combout  & ((\rfif.rdat2[16]~316_combout ))))) # (!Instr_IF_16 & (((\rfif.rdat2[16]~321_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[16]~323_combout ),
	.datac(\rfif.rdat2[16]~321_combout ),
	.datad(\rfif.rdat2[16]~316_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[16]~324_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[16]~324 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[16]~324 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N15
dffeas \regs[26][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][15] .is_wysiwyg = "true";
defparam \regs[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \rfif.rdat1[15]~320 (
// Equation(s):
// \rfif.rdat1[15]~320_combout  = (Instr_IF_24 & (((\regs[26][15]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[18][15]~q  & ((!Instr_IF_23))))

	.dataa(\regs[18][15]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[26][15]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~320_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~320 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[15]~320 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N27
dffeas \regs[30][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][15] .is_wysiwyg = "true";
defparam \regs[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N25
dffeas \regs[22][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][15] .is_wysiwyg = "true";
defparam \regs[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \rfif.rdat1[15]~321 (
// Equation(s):
// \rfif.rdat1[15]~321_combout  = (Instr_IF_23 & ((\rfif.rdat1[15]~320_combout  & (\regs[30][15]~q )) # (!\rfif.rdat1[15]~320_combout  & ((\regs[22][15]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[15]~320_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[15]~320_combout ),
	.datac(\regs[30][15]~q ),
	.datad(\regs[22][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~321_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~321 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[15]~321 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N29
dffeas \regs[20][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][15] .is_wysiwyg = "true";
defparam \regs[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N17
dffeas \regs[24][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][15] .is_wysiwyg = "true";
defparam \regs[24][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N11
dffeas \regs[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][15] .is_wysiwyg = "true";
defparam \regs[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[15]~324 (
// Equation(s):
// \rfif.rdat1[15]~324_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[24][15]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[16][15]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[24][15]~q ),
	.datad(\regs[16][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~324_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~324 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[15]~324 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[15]~325 (
// Equation(s):
// \rfif.rdat1[15]~325_combout  = (Instr_IF_23 & ((\rfif.rdat1[15]~324_combout  & (\regs[28][15]~q )) # (!\rfif.rdat1[15]~324_combout  & ((\regs[20][15]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[15]~324_combout ))))

	.dataa(\regs[28][15]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][15]~q ),
	.datad(\rfif.rdat1[15]~324_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~325_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~325 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[15]~325 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N17
dffeas \regs[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][15] .is_wysiwyg = "true";
defparam \regs[21][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N3
dffeas \regs[17][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][15] .is_wysiwyg = "true";
defparam \regs[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[15]~322 (
// Equation(s):
// \rfif.rdat1[15]~322_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][15]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & ((\regs[17][15]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[21][15]~q ),
	.datad(\regs[17][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~322_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~322 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[15]~322 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N29
dffeas \regs[25][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][15] .is_wysiwyg = "true";
defparam \regs[25][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N11
dffeas \regs[29][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][15] .is_wysiwyg = "true";
defparam \regs[29][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[15]~323 (
// Equation(s):
// \rfif.rdat1[15]~323_combout  = (Instr_IF_24 & ((\rfif.rdat1[15]~322_combout  & ((\regs[29][15]~q ))) # (!\rfif.rdat1[15]~322_combout  & (\regs[25][15]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[15]~322_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[15]~322_combout ),
	.datac(\regs[25][15]~q ),
	.datad(\regs[29][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~323_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~323 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[15]~323 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \rfif.rdat1[15]~326 (
// Equation(s):
// \rfif.rdat1[15]~326_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\rfif.rdat1[15]~323_combout ))) # (!Instr_IF_21 & (\rfif.rdat1[15]~325_combout ))))

	.dataa(\rfif.rdat1[15]~325_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[15]~323_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~326_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~326 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[15]~326 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N27
dffeas \regs[31][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][15] .is_wysiwyg = "true";
defparam \regs[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \regs[27][15]~feeder (
// Equation(s):
// \regs[27][15]~feeder_combout  = \input_b~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b15),
	.cin(gnd),
	.combout(\regs[27][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][15]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N9
dffeas \regs[27][15] (
	.clk(!CLK),
	.d(\regs[27][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][15] .is_wysiwyg = "true";
defparam \regs[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \regs[23][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][15] .is_wysiwyg = "true";
defparam \regs[23][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N13
dffeas \regs[19][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][15] .is_wysiwyg = "true";
defparam \regs[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[15]~327 (
// Equation(s):
// \rfif.rdat1[15]~327_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][15]~q )) # (!Instr_IF_23 & ((\regs[19][15]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][15]~q ),
	.datad(\regs[19][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~327_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~327 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[15]~327 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[15]~328 (
// Equation(s):
// \rfif.rdat1[15]~328_combout  = (\rfif.rdat1[15]~327_combout  & ((\regs[31][15]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[15]~327_combout  & (((\regs[27][15]~q  & Instr_IF_24))))

	.dataa(\regs[31][15]~q ),
	.datab(\regs[27][15]~q ),
	.datac(\rfif.rdat1[15]~327_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~328_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~328 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[15]~328 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N3
dffeas \regs[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][15] .is_wysiwyg = "true";
defparam \regs[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N19
dffeas \regs[11][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][15] .is_wysiwyg = "true";
defparam \regs[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N25
dffeas \regs[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][15] .is_wysiwyg = "true";
defparam \regs[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N29
dffeas \regs[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][15] .is_wysiwyg = "true";
defparam \regs[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[15]~330 (
// Equation(s):
// \rfif.rdat1[15]~330_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[9][15]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[8][15]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[9][15]~q ),
	.datad(\regs[8][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~330_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~330 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[15]~330 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \rfif.rdat1[15]~331 (
// Equation(s):
// \rfif.rdat1[15]~331_combout  = (Instr_IF_22 & ((\rfif.rdat1[15]~330_combout  & ((\regs[11][15]~q ))) # (!\rfif.rdat1[15]~330_combout  & (\regs[10][15]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[15]~330_combout ))))

	.dataa(\regs[10][15]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[11][15]~q ),
	.datad(\rfif.rdat1[15]~330_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~331_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~331 .lut_mask = 16'hF388;
defparam \rfif.rdat1[15]~331 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N15
dffeas \regs[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][15] .is_wysiwyg = "true";
defparam \regs[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N29
dffeas \regs[5][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][15] .is_wysiwyg = "true";
defparam \regs[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \rfif.rdat1[15]~333 (
// Equation(s):
// \rfif.rdat1[15]~333_combout  = (\rfif.rdat1[15]~332_combout  & ((\regs[7][15]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[15]~332_combout  & (((\regs[5][15]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[15]~332_combout ),
	.datab(\regs[7][15]~q ),
	.datac(\regs[5][15]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~333_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~333 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[15]~333 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N5
dffeas \regs[2][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][15] .is_wysiwyg = "true";
defparam \regs[2][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N9
dffeas \regs[3][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][15] .is_wysiwyg = "true";
defparam \regs[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N3
dffeas \regs[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][15] .is_wysiwyg = "true";
defparam \regs[1][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \regs[0][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][15] .is_wysiwyg = "true";
defparam \regs[0][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[15]~334 (
// Equation(s):
// \rfif.rdat1[15]~334_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][15]~q )) # (!Instr_IF_21 & ((\regs[0][15]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][15]~q ),
	.datad(\regs[0][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~334_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~334 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[15]~334 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[15]~335 (
// Equation(s):
// \rfif.rdat1[15]~335_combout  = (Instr_IF_22 & ((\rfif.rdat1[15]~334_combout  & ((\regs[3][15]~q ))) # (!\rfif.rdat1[15]~334_combout  & (\regs[2][15]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[15]~334_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[2][15]~q ),
	.datac(\regs[3][15]~q ),
	.datad(\rfif.rdat1[15]~334_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~335_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~335 .lut_mask = 16'hF588;
defparam \rfif.rdat1[15]~335 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[15]~336 (
// Equation(s):
// \rfif.rdat1[15]~336_combout  = (Instr_IF_23 & ((\rfif.rdat1[15]~333_combout ) # ((Instr_IF_24)))) # (!Instr_IF_23 & (((\rfif.rdat1[15]~335_combout  & !Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[15]~333_combout ),
	.datac(\rfif.rdat1[15]~335_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~336_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~336 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[15]~336 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N3
dffeas \regs[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][15] .is_wysiwyg = "true";
defparam \regs[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N29
dffeas \regs[14][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][15] .is_wysiwyg = "true";
defparam \regs[14][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[15]~337 (
// Equation(s):
// \rfif.rdat1[15]~337_combout  = (Instr_IF_22 & (((\regs[14][15]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[12][15]~q  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[12][15]~q ),
	.datac(\regs[14][15]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~337_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~337 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[15]~337 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N25
dffeas \regs[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][15] .is_wysiwyg = "true";
defparam \regs[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \regs[15][15]~feeder (
// Equation(s):
// \regs[15][15]~feeder_combout  = \input_b~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_b15),
	.cin(gnd),
	.combout(\regs[15][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][15]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N3
dffeas \regs[15][15] (
	.clk(!CLK),
	.d(\regs[15][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][15] .is_wysiwyg = "true";
defparam \regs[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \rfif.rdat1[15]~338 (
// Equation(s):
// \rfif.rdat1[15]~338_combout  = (\rfif.rdat1[15]~337_combout  & (((\regs[15][15]~q ) # (!Instr_IF_21)))) # (!\rfif.rdat1[15]~337_combout  & (\regs[13][15]~q  & ((Instr_IF_21))))

	.dataa(\rfif.rdat1[15]~337_combout ),
	.datab(\regs[13][15]~q ),
	.datac(\regs[15][15]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[15]~338_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[15]~338 .lut_mask = 16'hE4AA;
defparam \rfif.rdat1[15]~338 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[15]~346 (
// Equation(s):
// \rfif.rdat2[15]~346_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][15]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][15]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][15]~q ),
	.datad(\regs[9][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~346_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~346 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[15]~346 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[15]~347 (
// Equation(s):
// \rfif.rdat2[15]~347_combout  = (Instr_IF_17 & ((\rfif.rdat2[15]~346_combout  & ((\regs[11][15]~q ))) # (!\rfif.rdat2[15]~346_combout  & (\regs[10][15]~q )))) # (!Instr_IF_17 & (\rfif.rdat2[15]~346_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[15]~346_combout ),
	.datac(\regs[10][15]~q ),
	.datad(\regs[11][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~347_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~347 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[15]~347 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \rfif.rdat2[15]~353 (
// Equation(s):
// \rfif.rdat2[15]~353_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[14][15]~q ))) # (!Instr_IF_17 & (\regs[12][15]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][15]~q ),
	.datad(\regs[14][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~353_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~353 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[15]~353 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \rfif.rdat2[15]~354 (
// Equation(s):
// \rfif.rdat2[15]~354_combout  = (Instr_IF_16 & ((\rfif.rdat2[15]~353_combout  & ((\regs[15][15]~q ))) # (!\rfif.rdat2[15]~353_combout  & (\regs[13][15]~q )))) # (!Instr_IF_16 & (\rfif.rdat2[15]~353_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[15]~353_combout ),
	.datac(\regs[13][15]~q ),
	.datad(\regs[15][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~354_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~354 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[15]~354 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[15]~350 (
// Equation(s):
// \rfif.rdat2[15]~350_combout  = (Instr_IF_16 & ((\regs[1][15]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[0][15]~q  & !Instr_IF_17))))

	.dataa(\regs[1][15]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[0][15]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~350_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~350 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[15]~350 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \rfif.rdat2[15]~351 (
// Equation(s):
// \rfif.rdat2[15]~351_combout  = (Instr_IF_17 & ((\rfif.rdat2[15]~350_combout  & (\regs[3][15]~q )) # (!\rfif.rdat2[15]~350_combout  & ((\regs[2][15]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[15]~350_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[3][15]~q ),
	.datac(\regs[2][15]~q ),
	.datad(\rfif.rdat2[15]~350_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~351_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~351 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[15]~351 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N21
dffeas \regs[4][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][15] .is_wysiwyg = "true";
defparam \regs[4][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N3
dffeas \regs[6][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][15] .is_wysiwyg = "true";
defparam \regs[6][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \rfif.rdat2[15]~348 (
// Equation(s):
// \rfif.rdat2[15]~348_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][15]~q ))) # (!Instr_IF_17 & (\regs[4][15]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][15]~q ),
	.datad(\regs[6][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~348_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~348 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[15]~348 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \rfif.rdat2[15]~349 (
// Equation(s):
// \rfif.rdat2[15]~349_combout  = (Instr_IF_16 & ((\rfif.rdat2[15]~348_combout  & ((\regs[7][15]~q ))) # (!\rfif.rdat2[15]~348_combout  & (\regs[5][15]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[15]~348_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][15]~q ),
	.datac(\regs[7][15]~q ),
	.datad(\rfif.rdat2[15]~348_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~349_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~349 .lut_mask = 16'hF588;
defparam \rfif.rdat2[15]~349 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[15]~352 (
// Equation(s):
// \rfif.rdat2[15]~352_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\rfif.rdat2[15]~349_combout )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\rfif.rdat2[15]~351_combout )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[15]~351_combout ),
	.datad(\rfif.rdat2[15]~349_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~352_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~352 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[15]~352 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[15]~355 (
// Equation(s):
// \rfif.rdat2[15]~355_combout  = (Instr_IF_19 & ((\rfif.rdat2[15]~352_combout  & ((\rfif.rdat2[15]~354_combout ))) # (!\rfif.rdat2[15]~352_combout  & (\rfif.rdat2[15]~347_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[15]~352_combout ))))

	.dataa(\rfif.rdat2[15]~347_combout ),
	.datab(\rfif.rdat2[15]~354_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[15]~352_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~355_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~355 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[15]~355 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[15]~344 (
// Equation(s):
// \rfif.rdat2[15]~344_combout  = (\rfif.rdat2[15]~343_combout  & (((\regs[31][15]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[15]~343_combout  & (\regs[27][15]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[15]~343_combout ),
	.datab(\regs[27][15]~q ),
	.datac(\regs[31][15]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~344_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~344 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[15]~344 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N11
dffeas \regs[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][15] .is_wysiwyg = "true";
defparam \regs[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[15]~336 (
// Equation(s):
// \rfif.rdat2[15]~336_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[26][15]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & (\regs[18][15]~q )))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][15]~q ),
	.datad(\regs[26][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~336_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~336 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[15]~336 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \rfif.rdat2[15]~337 (
// Equation(s):
// \rfif.rdat2[15]~337_combout  = (Instr_IF_18 & ((\rfif.rdat2[15]~336_combout  & (\regs[30][15]~q )) # (!\rfif.rdat2[15]~336_combout  & ((\regs[22][15]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[15]~336_combout ))))

	.dataa(\regs[30][15]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][15]~q ),
	.datad(\rfif.rdat2[15]~336_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~337_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~337 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[15]~337 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \rfif.rdat2[15]~338 (
// Equation(s):
// \rfif.rdat2[15]~338_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][15]~q ))) # (!Instr_IF_18 & (\regs[17][15]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][15]~q ),
	.datad(\regs[21][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~338_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~338 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[15]~338 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[15]~339 (
// Equation(s):
// \rfif.rdat2[15]~339_combout  = (Instr_IF_19 & ((\rfif.rdat2[15]~338_combout  & ((\regs[29][15]~q ))) # (!\rfif.rdat2[15]~338_combout  & (\regs[25][15]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[15]~338_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][15]~q ),
	.datac(\regs[29][15]~q ),
	.datad(\rfif.rdat2[15]~338_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~339_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~339 .lut_mask = 16'hF588;
defparam \rfif.rdat2[15]~339 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N7
dffeas \regs[28][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][15] .is_wysiwyg = "true";
defparam \regs[28][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[15]~340 (
// Equation(s):
// \rfif.rdat2[15]~340_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][15]~q ))) # (!Instr_IF_19 & (\regs[16][15]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][15]~q ),
	.datad(\regs[24][15]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~340_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~340 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[15]~340 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[15]~341 (
// Equation(s):
// \rfif.rdat2[15]~341_combout  = (Instr_IF_18 & ((\rfif.rdat2[15]~340_combout  & ((\regs[28][15]~q ))) # (!\rfif.rdat2[15]~340_combout  & (\regs[20][15]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[15]~340_combout ))))

	.dataa(\regs[20][15]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][15]~q ),
	.datad(\rfif.rdat2[15]~340_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~341_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~341 .lut_mask = 16'hF388;
defparam \rfif.rdat2[15]~341 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N4
cycloneive_lcell_comb \rfif.rdat2[15]~342 (
// Equation(s):
// \rfif.rdat2[15]~342_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\rfif.rdat2[15]~339_combout )))) # (!Instr_IF_16 & (!Instr_IF_17 & ((\rfif.rdat2[15]~341_combout ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[15]~339_combout ),
	.datad(\rfif.rdat2[15]~341_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~342_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~342 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[15]~342 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[15]~345 (
// Equation(s):
// \rfif.rdat2[15]~345_combout  = (\rfif.rdat2[15]~342_combout  & ((\rfif.rdat2[15]~344_combout ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[15]~342_combout  & (((\rfif.rdat2[15]~337_combout  & Instr_IF_17))))

	.dataa(\rfif.rdat2[15]~344_combout ),
	.datab(\rfif.rdat2[15]~337_combout ),
	.datac(\rfif.rdat2[15]~342_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[15]~345_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[15]~345 .lut_mask = 16'hACF0;
defparam \rfif.rdat2[15]~345 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N23
dffeas \regs[17][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][14] .is_wysiwyg = "true";
defparam \regs[17][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N1
dffeas \regs[25][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][14] .is_wysiwyg = "true";
defparam \regs[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \rfif.rdat1[14]~340 (
// Equation(s):
// \rfif.rdat1[14]~340_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][14]~q ))) # (!Instr_IF_24 & (\regs[17][14]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[17][14]~q ),
	.datac(\regs[25][14]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~340_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~340 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[14]~340 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N15
dffeas \regs[29][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][14] .is_wysiwyg = "true";
defparam \regs[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N9
dffeas \regs[21][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][14] .is_wysiwyg = "true";
defparam \regs[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[14]~341 (
// Equation(s):
// \rfif.rdat1[14]~341_combout  = (Instr_IF_23 & ((\rfif.rdat1[14]~340_combout  & (\regs[29][14]~q )) # (!\rfif.rdat1[14]~340_combout  & ((\regs[21][14]~q ))))) # (!Instr_IF_23 & (\rfif.rdat1[14]~340_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[14]~340_combout ),
	.datac(\regs[29][14]~q ),
	.datad(\regs[21][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~341_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~341 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[14]~341 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N23
dffeas \regs[31][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][14] .is_wysiwyg = "true";
defparam \regs[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N9
dffeas \regs[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][14] .is_wysiwyg = "true";
defparam \regs[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N11
dffeas \regs[27][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][14] .is_wysiwyg = "true";
defparam \regs[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N7
dffeas \regs[19][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][14] .is_wysiwyg = "true";
defparam \regs[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[14]~347 (
// Equation(s):
// \rfif.rdat1[14]~347_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][14]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][14]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][14]~q ),
	.datad(\regs[19][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~347_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~347 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[14]~347 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N8
cycloneive_lcell_comb \rfif.rdat1[14]~348 (
// Equation(s):
// \rfif.rdat1[14]~348_combout  = (Instr_IF_23 & ((\rfif.rdat1[14]~347_combout  & (\regs[31][14]~q )) # (!\rfif.rdat1[14]~347_combout  & ((\regs[23][14]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[14]~347_combout ))))

	.dataa(\regs[31][14]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[23][14]~q ),
	.datad(\rfif.rdat1[14]~347_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~348_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~348 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[14]~348 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N17
dffeas \regs[24][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][14] .is_wysiwyg = "true";
defparam \regs[24][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N15
dffeas \regs[28][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][14] .is_wysiwyg = "true";
defparam \regs[28][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[14]~345 (
// Equation(s):
// \rfif.rdat1[14]~345_combout  = (\rfif.rdat1[14]~344_combout  & (((\regs[28][14]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[14]~344_combout  & (Instr_IF_24 & (\regs[24][14]~q )))

	.dataa(\rfif.rdat1[14]~344_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[24][14]~q ),
	.datad(\regs[28][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~345_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~345 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[14]~345 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N15
dffeas \regs[30][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][14] .is_wysiwyg = "true";
defparam \regs[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \regs[26][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][14] .is_wysiwyg = "true";
defparam \regs[26][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N3
dffeas \regs[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][14] .is_wysiwyg = "true";
defparam \regs[18][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N29
dffeas \regs[22][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][14] .is_wysiwyg = "true";
defparam \regs[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \rfif.rdat1[14]~342 (
// Equation(s):
// \rfif.rdat1[14]~342_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][14]~q ))) # (!Instr_IF_23 & (\regs[18][14]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[18][14]~q ),
	.datac(\regs[22][14]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~342_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~342 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[14]~342 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \rfif.rdat1[14]~343 (
// Equation(s):
// \rfif.rdat1[14]~343_combout  = (Instr_IF_24 & ((\rfif.rdat1[14]~342_combout  & (\regs[30][14]~q )) # (!\rfif.rdat1[14]~342_combout  & ((\regs[26][14]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[14]~342_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[30][14]~q ),
	.datac(\regs[26][14]~q ),
	.datad(\rfif.rdat1[14]~342_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~343_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~343 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[14]~343 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[14]~346 (
// Equation(s):
// \rfif.rdat1[14]~346_combout  = (Instr_IF_22 & (((\rfif.rdat1[14]~343_combout ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\rfif.rdat1[14]~345_combout  & ((!Instr_IF_21))))

	.dataa(\rfif.rdat1[14]~345_combout ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[14]~343_combout ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~346_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~346 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[14]~346 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N25
dffeas \regs[13][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][14] .is_wysiwyg = "true";
defparam \regs[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \rfif.rdat1[14]~357 (
// Equation(s):
// \rfif.rdat1[14]~357_combout  = (Instr_IF_21 & (((\regs[13][14]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][14]~q  & ((!Instr_IF_22))))

	.dataa(\regs[12][14]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][14]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~357_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~357 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[14]~357 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N11
dffeas \regs[14][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][14] .is_wysiwyg = "true";
defparam \regs[14][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N9
dffeas \regs[15][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][14] .is_wysiwyg = "true";
defparam \regs[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[14]~358 (
// Equation(s):
// \rfif.rdat1[14]~358_combout  = (Instr_IF_22 & ((\rfif.rdat1[14]~357_combout  & ((\regs[15][14]~q ))) # (!\rfif.rdat1[14]~357_combout  & (\regs[14][14]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[14]~357_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[14]~357_combout ),
	.datac(\regs[14][14]~q ),
	.datad(\regs[15][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~358_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~358 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[14]~358 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N23
dffeas \regs[7][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][14] .is_wysiwyg = "true";
defparam \regs[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N15
dffeas \regs[6][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][14] .is_wysiwyg = "true";
defparam \regs[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N17
dffeas \regs[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][14] .is_wysiwyg = "true";
defparam \regs[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[14]~350 (
// Equation(s):
// \rfif.rdat1[14]~350_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[5][14]~q )) # (!Instr_IF_21 & ((\regs[4][14]~q )))))

	.dataa(\regs[5][14]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[4][14]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~350_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~350 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[14]~350 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[14]~351 (
// Equation(s):
// \rfif.rdat1[14]~351_combout  = (Instr_IF_22 & ((\rfif.rdat1[14]~350_combout  & (\regs[7][14]~q )) # (!\rfif.rdat1[14]~350_combout  & ((\regs[6][14]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[14]~350_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[7][14]~q ),
	.datac(\regs[6][14]~q ),
	.datad(\rfif.rdat1[14]~350_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~351_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~351 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[14]~351 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \regs[11][14]~feeder (
// Equation(s):
// \regs[11][14]~feeder_combout  = \input_b~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b16),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][14]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N3
dffeas \regs[11][14] (
	.clk(!CLK),
	.d(\regs[11][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][14] .is_wysiwyg = "true";
defparam \regs[11][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \regs[9][14]~feeder (
// Equation(s):
// \regs[9][14]~feeder_combout  = \input_b~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b16),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][14]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N5
dffeas \regs[9][14] (
	.clk(!CLK),
	.d(\regs[9][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][14] .is_wysiwyg = "true";
defparam \regs[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N5
dffeas \regs[8][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][14] .is_wysiwyg = "true";
defparam \regs[8][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N19
dffeas \regs[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][14] .is_wysiwyg = "true";
defparam \regs[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \rfif.rdat1[14]~352 (
// Equation(s):
// \rfif.rdat1[14]~352_combout  = (Instr_IF_22 & (((\regs[10][14]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[8][14]~q  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[8][14]~q ),
	.datac(\regs[10][14]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~352_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~352 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[14]~352 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \rfif.rdat1[14]~353 (
// Equation(s):
// \rfif.rdat1[14]~353_combout  = (Instr_IF_21 & ((\rfif.rdat1[14]~352_combout  & (\regs[11][14]~q )) # (!\rfif.rdat1[14]~352_combout  & ((\regs[9][14]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[14]~352_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][14]~q ),
	.datac(\regs[9][14]~q ),
	.datad(\rfif.rdat1[14]~352_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~353_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~353 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[14]~353 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N5
dffeas \regs[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][14] .is_wysiwyg = "true";
defparam \regs[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N1
dffeas \regs[2][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][14] .is_wysiwyg = "true";
defparam \regs[2][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[14]~354 (
// Equation(s):
// \rfif.rdat1[14]~354_combout  = (Instr_IF_22 & (((\regs[2][14]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[0][14]~q  & ((!Instr_IF_21))))

	.dataa(\regs[0][14]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[2][14]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~354_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~354 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[14]~354 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[14]~355 (
// Equation(s):
// \rfif.rdat1[14]~355_combout  = (Instr_IF_21 & ((\rfif.rdat1[14]~354_combout  & (\regs[3][14]~q )) # (!\rfif.rdat1[14]~354_combout  & ((\regs[1][14]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[14]~354_combout ))))

	.dataa(\regs[3][14]~q ),
	.datab(\regs[1][14]~q ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[14]~354_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~355_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~355 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[14]~355 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[14]~356 (
// Equation(s):
// \rfif.rdat1[14]~356_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\rfif.rdat1[14]~353_combout )) # (!Instr_IF_24 & ((\rfif.rdat1[14]~355_combout )))))

	.dataa(\rfif.rdat1[14]~353_combout ),
	.datab(Instr_IF_23),
	.datac(\rfif.rdat1[14]~355_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[14]~356_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[14]~356 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[14]~356 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N8
cycloneive_lcell_comb \rfif.rdat2[14]~358 (
// Equation(s):
// \rfif.rdat2[14]~358_combout  = (\rfif.rdat2[14]~357_combout  & (((\regs[29][14]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[14]~357_combout  & (Instr_IF_18 & (\regs[21][14]~q )))

	.dataa(\rfif.rdat2[14]~357_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[21][14]~q ),
	.datad(\regs[29][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~358_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~358 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[14]~358 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N17
dffeas \regs[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][14] .is_wysiwyg = "true";
defparam \regs[20][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[14]~361 (
// Equation(s):
// \rfif.rdat2[14]~361_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[20][14]~q ))) # (!Instr_IF_18 & (\regs[16][14]~q ))))

	.dataa(\regs[16][14]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[20][14]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~361_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~361 .lut_mask = 16'hFC22;
defparam \rfif.rdat2[14]~361 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[14]~362 (
// Equation(s):
// \rfif.rdat2[14]~362_combout  = (Instr_IF_19 & ((\rfif.rdat2[14]~361_combout  & ((\regs[28][14]~q ))) # (!\rfif.rdat2[14]~361_combout  & (\regs[24][14]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[14]~361_combout ))))

	.dataa(\regs[24][14]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[28][14]~q ),
	.datad(\rfif.rdat2[14]~361_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~362_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~362 .lut_mask = 16'hF388;
defparam \rfif.rdat2[14]~362 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \rfif.rdat2[14]~359 (
// Equation(s):
// \rfif.rdat2[14]~359_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][14]~q ))) # (!Instr_IF_18 & (\regs[18][14]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][14]~q ),
	.datad(\regs[22][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~359_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~359 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[14]~359 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[14]~360 (
// Equation(s):
// \rfif.rdat2[14]~360_combout  = (Instr_IF_19 & ((\rfif.rdat2[14]~359_combout  & ((\regs[30][14]~q ))) # (!\rfif.rdat2[14]~359_combout  & (\regs[26][14]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[14]~359_combout ))))

	.dataa(\regs[26][14]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[30][14]~q ),
	.datad(\rfif.rdat2[14]~359_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~360_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~360 .lut_mask = 16'hF388;
defparam \rfif.rdat2[14]~360 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[14]~363 (
// Equation(s):
// \rfif.rdat2[14]~363_combout  = (Instr_IF_17 & (((\rfif.rdat2[14]~360_combout ) # (Instr_IF_16)))) # (!Instr_IF_17 & (\rfif.rdat2[14]~362_combout  & ((!Instr_IF_16))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[14]~362_combout ),
	.datac(\rfif.rdat2[14]~360_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~363_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~363 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[14]~363 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[14]~364 (
// Equation(s):
// \rfif.rdat2[14]~364_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[27][14]~q ))) # (!Instr_IF_19 & (\regs[19][14]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][14]~q ),
	.datad(\regs[27][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~364_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~364 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[14]~364 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[14]~365 (
// Equation(s):
// \rfif.rdat2[14]~365_combout  = (Instr_IF_18 & ((\rfif.rdat2[14]~364_combout  & ((\regs[31][14]~q ))) # (!\rfif.rdat2[14]~364_combout  & (\regs[23][14]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[14]~364_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][14]~q ),
	.datac(\regs[31][14]~q ),
	.datad(\rfif.rdat2[14]~364_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~365_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~365 .lut_mask = 16'hF588;
defparam \rfif.rdat2[14]~365 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[14]~366 (
// Equation(s):
// \rfif.rdat2[14]~366_combout  = (Instr_IF_16 & ((\rfif.rdat2[14]~363_combout  & ((\rfif.rdat2[14]~365_combout ))) # (!\rfif.rdat2[14]~363_combout  & (\rfif.rdat2[14]~358_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[14]~363_combout ))))

	.dataa(\rfif.rdat2[14]~358_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[14]~363_combout ),
	.datad(\rfif.rdat2[14]~365_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~366_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~366 .lut_mask = 16'hF838;
defparam \rfif.rdat2[14]~366 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N1
dffeas \regs[5][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][14] .is_wysiwyg = "true";
defparam \regs[5][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[14]~367 (
// Equation(s):
// \rfif.rdat2[14]~367_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[5][14]~q )) # (!Instr_IF_16 & ((\regs[4][14]~q )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[5][14]~q ),
	.datad(\regs[4][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~367_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~367 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[14]~367 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[14]~368 (
// Equation(s):
// \rfif.rdat2[14]~368_combout  = (Instr_IF_17 & ((\rfif.rdat2[14]~367_combout  & ((\regs[7][14]~q ))) # (!\rfif.rdat2[14]~367_combout  & (\regs[6][14]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[14]~367_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[6][14]~q ),
	.datac(\regs[7][14]~q ),
	.datad(\rfif.rdat2[14]~367_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~368_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~368 .lut_mask = 16'hF588;
defparam \rfif.rdat2[14]~368 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N23
dffeas \regs[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][14] .is_wysiwyg = "true";
defparam \regs[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \rfif.rdat2[14]~374 (
// Equation(s):
// \rfif.rdat2[14]~374_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][14]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][14]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][14]~q ),
	.datad(\regs[13][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~374_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~374 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[14]~374 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[14]~375 (
// Equation(s):
// \rfif.rdat2[14]~375_combout  = (Instr_IF_17 & ((\rfif.rdat2[14]~374_combout  & (\regs[15][14]~q )) # (!\rfif.rdat2[14]~374_combout  & ((\regs[14][14]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[14]~374_combout ))))

	.dataa(\regs[15][14]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[14][14]~q ),
	.datad(\rfif.rdat2[14]~374_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~375_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~375 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[14]~375 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \rfif.rdat2[14]~369 (
// Equation(s):
// \rfif.rdat2[14]~369_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[10][14]~q )) # (!Instr_IF_17 & ((\regs[8][14]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[10][14]~q ),
	.datac(\regs[8][14]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~369_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~369 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[14]~369 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[14]~370 (
// Equation(s):
// \rfif.rdat2[14]~370_combout  = (Instr_IF_16 & ((\rfif.rdat2[14]~369_combout  & ((\regs[11][14]~q ))) # (!\rfif.rdat2[14]~369_combout  & (\regs[9][14]~q )))) # (!Instr_IF_16 & (\rfif.rdat2[14]~369_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[14]~369_combout ),
	.datac(\regs[9][14]~q ),
	.datad(\regs[11][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~370_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~370 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[14]~370 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \regs[0][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_b16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][14] .is_wysiwyg = "true";
defparam \regs[0][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[14]~371 (
// Equation(s):
// \rfif.rdat2[14]~371_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][14]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][14]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][14]~q ),
	.datad(\regs[2][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~371_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~371 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[14]~371 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \regs[3][14]~feeder (
// Equation(s):
// \regs[3][14]~feeder_combout  = \input_b~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_b16),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][14]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N11
dffeas \regs[3][14] (
	.clk(!CLK),
	.d(\regs[3][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][14] .is_wysiwyg = "true";
defparam \regs[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[14]~372 (
// Equation(s):
// \rfif.rdat2[14]~372_combout  = (Instr_IF_16 & ((\rfif.rdat2[14]~371_combout  & ((\regs[3][14]~q ))) # (!\rfif.rdat2[14]~371_combout  & (\regs[1][14]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[14]~371_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][14]~q ),
	.datac(\rfif.rdat2[14]~371_combout ),
	.datad(\regs[3][14]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~372_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~372 .lut_mask = 16'hF858;
defparam \rfif.rdat2[14]~372 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[14]~373 (
// Equation(s):
// \rfif.rdat2[14]~373_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\rfif.rdat2[14]~370_combout )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\rfif.rdat2[14]~372_combout ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[14]~370_combout ),
	.datad(\rfif.rdat2[14]~372_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~373_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~373 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[14]~373 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[14]~376 (
// Equation(s):
// \rfif.rdat2[14]~376_combout  = (Instr_IF_18 & ((\rfif.rdat2[14]~373_combout  & ((\rfif.rdat2[14]~375_combout ))) # (!\rfif.rdat2[14]~373_combout  & (\rfif.rdat2[14]~368_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[14]~373_combout ))))

	.dataa(\rfif.rdat2[14]~368_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[14]~375_combout ),
	.datad(\rfif.rdat2[14]~373_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[14]~376_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[14]~376 .lut_mask = 16'hF388;
defparam \rfif.rdat2[14]~376 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N19
dffeas \regs[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][13] .is_wysiwyg = "true";
defparam \regs[18][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N21
dffeas \regs[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][13] .is_wysiwyg = "true";
defparam \regs[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \rfif.rdat2[13]~378 (
// Equation(s):
// \rfif.rdat2[13]~378_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[26][13]~q ))) # (!Instr_IF_19 & (\regs[18][13]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[18][13]~q ),
	.datac(\regs[26][13]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~378_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~378 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[13]~378 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N5
dffeas \regs[22][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][13] .is_wysiwyg = "true";
defparam \regs[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N31
dffeas \regs[30][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][13] .is_wysiwyg = "true";
defparam \regs[30][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[13]~379 (
// Equation(s):
// \rfif.rdat2[13]~379_combout  = (Instr_IF_18 & ((\rfif.rdat2[13]~378_combout  & ((\regs[30][13]~q ))) # (!\rfif.rdat2[13]~378_combout  & (\regs[22][13]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[13]~378_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[13]~378_combout ),
	.datac(\regs[22][13]~q ),
	.datad(\regs[30][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~379_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~379 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[13]~379 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N25
dffeas \regs[25][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][13] .is_wysiwyg = "true";
defparam \regs[25][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N3
dffeas \regs[29][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][13] .is_wysiwyg = "true";
defparam \regs[29][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N27
dffeas \regs[17][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][13] .is_wysiwyg = "true";
defparam \regs[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N0
cycloneive_lcell_comb \regs[21][13]~feeder (
// Equation(s):
// \regs[21][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[21][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[21][13]~feeder .lut_mask = 16'hF0F0;
defparam \regs[21][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N1
dffeas \regs[21][13] (
	.clk(!CLK),
	.d(\regs[21][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][13] .is_wysiwyg = "true";
defparam \regs[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[13]~380 (
// Equation(s):
// \rfif.rdat2[13]~380_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[21][13]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[17][13]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[17][13]~q ),
	.datad(\regs[21][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~380_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~380 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[13]~380 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[13]~381 (
// Equation(s):
// \rfif.rdat2[13]~381_combout  = (Instr_IF_19 & ((\rfif.rdat2[13]~380_combout  & ((\regs[29][13]~q ))) # (!\rfif.rdat2[13]~380_combout  & (\regs[25][13]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[13]~380_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][13]~q ),
	.datac(\regs[29][13]~q ),
	.datad(\rfif.rdat2[13]~380_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~381_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~381 .lut_mask = 16'hF588;
defparam \rfif.rdat2[13]~381 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[13]~384 (
// Equation(s):
// \rfif.rdat2[13]~384_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\rfif.rdat2[13]~381_combout ))) # (!Instr_IF_16 & (\rfif.rdat2[13]~383_combout ))))

	.dataa(\rfif.rdat2[13]~383_combout ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[13]~381_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~384_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~384 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[13]~384 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N14
cycloneive_lcell_comb \regs[27][13]~feeder (
// Equation(s):
// \regs[27][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[27][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N15
dffeas \regs[27][13] (
	.clk(!CLK),
	.d(\regs[27][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][13] .is_wysiwyg = "true";
defparam \regs[27][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N8
cycloneive_lcell_comb \regs[23][13]~feeder (
// Equation(s):
// \regs[23][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[23][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[23][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[23][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N9
dffeas \regs[23][13] (
	.clk(!CLK),
	.d(\regs[23][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][13] .is_wysiwyg = "true";
defparam \regs[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N25
dffeas \regs[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][13] .is_wysiwyg = "true";
defparam \regs[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \rfif.rdat2[13]~385 (
// Equation(s):
// \rfif.rdat2[13]~385_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[23][13]~q )) # (!Instr_IF_18 & ((\regs[19][13]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[23][13]~q ),
	.datac(\regs[19][13]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~385_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~385 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[13]~385 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \rfif.rdat2[13]~386 (
// Equation(s):
// \rfif.rdat2[13]~386_combout  = (Instr_IF_19 & ((\rfif.rdat2[13]~385_combout  & (\regs[31][13]~q )) # (!\rfif.rdat2[13]~385_combout  & ((\regs[27][13]~q ))))) # (!Instr_IF_19 & (((\rfif.rdat2[13]~385_combout ))))

	.dataa(\regs[31][13]~q ),
	.datab(\regs[27][13]~q ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[13]~385_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~386_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~386 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[13]~386 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[13]~387 (
// Equation(s):
// \rfif.rdat2[13]~387_combout  = (Instr_IF_17 & ((\rfif.rdat2[13]~384_combout  & ((\rfif.rdat2[13]~386_combout ))) # (!\rfif.rdat2[13]~384_combout  & (\rfif.rdat2[13]~379_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[13]~384_combout ))))

	.dataa(\rfif.rdat2[13]~379_combout ),
	.datab(Instr_IF_17),
	.datac(\rfif.rdat2[13]~384_combout ),
	.datad(\rfif.rdat2[13]~386_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~387_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~387 .lut_mask = 16'hF838;
defparam \rfif.rdat2[13]~387 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \regs[2][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][13] .is_wysiwyg = "true";
defparam \regs[2][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N11
dffeas \regs[0][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][13] .is_wysiwyg = "true";
defparam \regs[0][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \regs[1][13]~feeder (
// Equation(s):
// \regs[1][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[1][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[1][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N25
dffeas \regs[1][13] (
	.clk(!CLK),
	.d(\regs[1][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][13] .is_wysiwyg = "true";
defparam \regs[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[13]~392 (
// Equation(s):
// \rfif.rdat2[13]~392_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][13]~q ))) # (!Instr_IF_16 & (\regs[0][13]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][13]~q ),
	.datad(\regs[1][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~392_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~392 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[13]~392 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \rfif.rdat2[13]~393 (
// Equation(s):
// \rfif.rdat2[13]~393_combout  = (Instr_IF_17 & ((\rfif.rdat2[13]~392_combout  & (\regs[3][13]~q )) # (!\rfif.rdat2[13]~392_combout  & ((\regs[2][13]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[13]~392_combout ))))

	.dataa(\regs[3][13]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[2][13]~q ),
	.datad(\rfif.rdat2[13]~392_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~393_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~393 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[13]~393 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[13]~394 (
// Equation(s):
// \rfif.rdat2[13]~394_combout  = (Instr_IF_18 & ((\rfif.rdat2[13]~391_combout ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((!Instr_IF_19 & \rfif.rdat2[13]~393_combout ))))

	.dataa(\rfif.rdat2[13]~391_combout ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[13]~393_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~394_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~394 .lut_mask = 16'hCBC8;
defparam \rfif.rdat2[13]~394 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N7
dffeas \regs[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][13] .is_wysiwyg = "true";
defparam \regs[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \regs[15][13]~feeder (
// Equation(s):
// \regs[15][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N31
dffeas \regs[15][13] (
	.clk(!CLK),
	.d(\regs[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][13] .is_wysiwyg = "true";
defparam \regs[15][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N29
dffeas \regs[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][13] .is_wysiwyg = "true";
defparam \regs[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \regs[14][13]~feeder (
// Equation(s):
// \regs[14][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[14][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N29
dffeas \regs[14][13] (
	.clk(!CLK),
	.d(\regs[14][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][13] .is_wysiwyg = "true";
defparam \regs[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[13]~395 (
// Equation(s):
// \rfif.rdat2[13]~395_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][13]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][13]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][13]~q ),
	.datad(\regs[14][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~395_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~395 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[13]~395 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[13]~396 (
// Equation(s):
// \rfif.rdat2[13]~396_combout  = (Instr_IF_16 & ((\rfif.rdat2[13]~395_combout  & ((\regs[15][13]~q ))) # (!\rfif.rdat2[13]~395_combout  & (\regs[13][13]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[13]~395_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[13][13]~q ),
	.datac(\regs[15][13]~q ),
	.datad(\rfif.rdat2[13]~395_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~396_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~396 .lut_mask = 16'hF588;
defparam \rfif.rdat2[13]~396 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N27
dffeas \regs[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][13] .is_wysiwyg = "true";
defparam \regs[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N14
cycloneive_lcell_comb \regs[11][13]~feeder (
// Equation(s):
// \regs[11][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[11][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[11][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N15
dffeas \regs[11][13] (
	.clk(!CLK),
	.d(\regs[11][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][13] .is_wysiwyg = "true";
defparam \regs[11][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N1
dffeas \regs[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][13] .is_wysiwyg = "true";
defparam \regs[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N16
cycloneive_lcell_comb \regs[9][13]~feeder (
// Equation(s):
// \regs[9][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[9][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N17
dffeas \regs[9][13] (
	.clk(!CLK),
	.d(\regs[9][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][13] .is_wysiwyg = "true";
defparam \regs[9][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[13]~388 (
// Equation(s):
// \rfif.rdat2[13]~388_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][13]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][13]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][13]~q ),
	.datad(\regs[9][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~388_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~388 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[13]~388 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N12
cycloneive_lcell_comb \rfif.rdat2[13]~389 (
// Equation(s):
// \rfif.rdat2[13]~389_combout  = (Instr_IF_17 & ((\rfif.rdat2[13]~388_combout  & ((\regs[11][13]~q ))) # (!\rfif.rdat2[13]~388_combout  & (\regs[10][13]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[13]~388_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[10][13]~q ),
	.datac(\regs[11][13]~q ),
	.datad(\rfif.rdat2[13]~388_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~389_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~389 .lut_mask = 16'hF588;
defparam \rfif.rdat2[13]~389 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[13]~397 (
// Equation(s):
// \rfif.rdat2[13]~397_combout  = (\rfif.rdat2[13]~394_combout  & ((\rfif.rdat2[13]~396_combout ) # ((!Instr_IF_19)))) # (!\rfif.rdat2[13]~394_combout  & (((Instr_IF_19 & \rfif.rdat2[13]~389_combout ))))

	.dataa(\rfif.rdat2[13]~394_combout ),
	.datab(\rfif.rdat2[13]~396_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[13]~389_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[13]~397_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[13]~397 .lut_mask = 16'hDA8A;
defparam \rfif.rdat2[13]~397 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \rfif.rdat1[13]~362 (
// Equation(s):
// \rfif.rdat1[13]~362_combout  = (Instr_IF_23 & ((\regs[22][13]~q ) # ((Instr_IF_24)))) # (!Instr_IF_23 & (((\regs[18][13]~q  & !Instr_IF_24))))

	.dataa(\regs[22][13]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[18][13]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~362_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~362 .lut_mask = 16'hCCB8;
defparam \rfif.rdat1[13]~362 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \rfif.rdat1[13]~363 (
// Equation(s):
// \rfif.rdat1[13]~363_combout  = (Instr_IF_24 & ((\rfif.rdat1[13]~362_combout  & ((\regs[30][13]~q ))) # (!\rfif.rdat1[13]~362_combout  & (\regs[26][13]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[13]~362_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[26][13]~q ),
	.datac(\regs[30][13]~q ),
	.datad(\rfif.rdat1[13]~362_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~363_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~363 .lut_mask = 16'hF588;
defparam \rfif.rdat1[13]~363 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N31
dffeas \regs[28][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][13] .is_wysiwyg = "true";
defparam \regs[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N21
dffeas \regs[24][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][13] .is_wysiwyg = "true";
defparam \regs[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[13]~365 (
// Equation(s):
// \rfif.rdat1[13]~365_combout  = (\rfif.rdat1[13]~364_combout  & ((\regs[28][13]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[13]~364_combout  & (((\regs[24][13]~q  & Instr_IF_24))))

	.dataa(\rfif.rdat1[13]~364_combout ),
	.datab(\regs[28][13]~q ),
	.datac(\regs[24][13]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~365_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~365 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[13]~365 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N30
cycloneive_lcell_comb \rfif.rdat1[13]~366 (
// Equation(s):
// \rfif.rdat1[13]~366_combout  = (Instr_IF_22 & ((\rfif.rdat1[13]~363_combout ) # ((Instr_IF_21)))) # (!Instr_IF_22 & (((!Instr_IF_21 & \rfif.rdat1[13]~365_combout ))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[13]~363_combout ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[13]~365_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~366_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~366 .lut_mask = 16'hADA8;
defparam \rfif.rdat1[13]~366 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[13]~360 (
// Equation(s):
// \rfif.rdat1[13]~360_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][13]~q ))) # (!Instr_IF_24 & (\regs[17][13]~q ))))

	.dataa(\regs[17][13]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[25][13]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~360_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~360 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[13]~360 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \rfif.rdat1[13]~361 (
// Equation(s):
// \rfif.rdat1[13]~361_combout  = (Instr_IF_23 & ((\rfif.rdat1[13]~360_combout  & ((\regs[29][13]~q ))) # (!\rfif.rdat1[13]~360_combout  & (\regs[21][13]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[13]~360_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[21][13]~q ),
	.datac(\regs[29][13]~q ),
	.datad(\rfif.rdat1[13]~360_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~361_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~361 .lut_mask = 16'hF588;
defparam \rfif.rdat1[13]~361 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N10
cycloneive_lcell_comb \rfif.rdat1[13]~367 (
// Equation(s):
// \rfif.rdat1[13]~367_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[27][13]~q )) # (!Instr_IF_24 & ((\regs[19][13]~q )))))

	.dataa(Instr_IF_23),
	.datab(\regs[27][13]~q ),
	.datac(\regs[19][13]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~367_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~367 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[13]~367 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \regs[31][13]~feeder (
// Equation(s):
// \regs[31][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a1),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][13]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N31
dffeas \regs[31][13] (
	.clk(!CLK),
	.d(\regs[31][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][13] .is_wysiwyg = "true";
defparam \regs[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[13]~368 (
// Equation(s):
// \rfif.rdat1[13]~368_combout  = (\rfif.rdat1[13]~367_combout  & (((\regs[31][13]~q ) # (!Instr_IF_23)))) # (!\rfif.rdat1[13]~367_combout  & (\regs[23][13]~q  & ((Instr_IF_23))))

	.dataa(\rfif.rdat1[13]~367_combout ),
	.datab(\regs[23][13]~q ),
	.datac(\regs[31][13]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~368_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~368 .lut_mask = 16'hE4AA;
defparam \rfif.rdat1[13]~368 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \regs[7][13]~feeder (
// Equation(s):
// \regs[7][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[7][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[7][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N9
dffeas \regs[7][13] (
	.clk(!CLK),
	.d(\regs[7][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][13] .is_wysiwyg = "true";
defparam \regs[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N23
dffeas \regs[6][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][13] .is_wysiwyg = "true";
defparam \regs[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N19
dffeas \regs[5][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][13] .is_wysiwyg = "true";
defparam \regs[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[13]~370 (
// Equation(s):
// \rfif.rdat1[13]~370_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][13]~q ))) # (!Instr_IF_21 & (\regs[4][13]~q ))))

	.dataa(\regs[4][13]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[5][13]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~370_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~370 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[13]~370 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \rfif.rdat1[13]~371 (
// Equation(s):
// \rfif.rdat1[13]~371_combout  = (Instr_IF_22 & ((\rfif.rdat1[13]~370_combout  & (\regs[7][13]~q )) # (!\rfif.rdat1[13]~370_combout  & ((\regs[6][13]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[13]~370_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[7][13]~q ),
	.datac(\regs[6][13]~q ),
	.datad(\rfif.rdat1[13]~370_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~371_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~371 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[13]~371 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[13]~377 (
// Equation(s):
// \rfif.rdat1[13]~377_combout  = (Instr_IF_21 & (((\regs[13][13]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][13]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][13]~q ),
	.datac(\regs[13][13]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~377_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~377 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[13]~377 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[13]~378 (
// Equation(s):
// \rfif.rdat1[13]~378_combout  = (Instr_IF_22 & ((\rfif.rdat1[13]~377_combout  & (\regs[15][13]~q )) # (!\rfif.rdat1[13]~377_combout  & ((\regs[14][13]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[13]~377_combout ))))

	.dataa(\regs[15][13]~q ),
	.datab(\regs[14][13]~q ),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[13]~377_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~378_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~378 .lut_mask = 16'hAFC0;
defparam \rfif.rdat1[13]~378 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[13]~374 (
// Equation(s):
// \rfif.rdat1[13]~374_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][13]~q )) # (!Instr_IF_22 & ((\regs[0][13]~q )))))

	.dataa(Instr_IF_21),
	.datab(\regs[2][13]~q ),
	.datac(\regs[0][13]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~374_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~374 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[13]~374 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \regs[3][13]~feeder (
// Equation(s):
// \regs[3][13]~feeder_combout  = \input_a~96_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a1),
	.cin(gnd),
	.combout(\regs[3][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][13]~feeder .lut_mask = 16'hFF00;
defparam \regs[3][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N15
dffeas \regs[3][13] (
	.clk(!CLK),
	.d(\regs[3][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][13] .is_wysiwyg = "true";
defparam \regs[3][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \rfif.rdat1[13]~375 (
// Equation(s):
// \rfif.rdat1[13]~375_combout  = (Instr_IF_21 & ((\rfif.rdat1[13]~374_combout  & (\regs[3][13]~q )) # (!\rfif.rdat1[13]~374_combout  & ((\regs[1][13]~q ))))) # (!Instr_IF_21 & (\rfif.rdat1[13]~374_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[13]~374_combout ),
	.datac(\regs[3][13]~q ),
	.datad(\regs[1][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~375_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~375 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[13]~375 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \rfif.rdat1[13]~372 (
// Equation(s):
// \rfif.rdat1[13]~372_combout  = (Instr_IF_22 & (((\regs[10][13]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[8][13]~q  & ((!Instr_IF_21))))

	.dataa(\regs[8][13]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[10][13]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~372_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~372 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[13]~372 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[13]~373 (
// Equation(s):
// \rfif.rdat1[13]~373_combout  = (Instr_IF_21 & ((\rfif.rdat1[13]~372_combout  & ((\regs[11][13]~q ))) # (!\rfif.rdat1[13]~372_combout  & (\regs[9][13]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[13]~372_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[9][13]~q ),
	.datac(\rfif.rdat1[13]~372_combout ),
	.datad(\regs[11][13]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~373_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~373 .lut_mask = 16'hF858;
defparam \rfif.rdat1[13]~373 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[13]~376 (
// Equation(s):
// \rfif.rdat1[13]~376_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[13]~373_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[13]~375_combout ))))

	.dataa(\rfif.rdat1[13]~375_combout ),
	.datab(Instr_IF_23),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[13]~373_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[13]~376_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[13]~376 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[13]~376 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N21
dffeas \regs[21][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][12] .is_wysiwyg = "true";
defparam \regs[21][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N9
dffeas \regs[25][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][12] .is_wysiwyg = "true";
defparam \regs[25][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \rfif.rdat2[12]~399 (
// Equation(s):
// \rfif.rdat2[12]~399_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][12]~q ))) # (!Instr_IF_19 & (\regs[17][12]~q ))))

	.dataa(\regs[17][12]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[25][12]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~399_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~399 .lut_mask = 16'hFC22;
defparam \rfif.rdat2[12]~399 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[12]~400 (
// Equation(s):
// \rfif.rdat2[12]~400_combout  = (Instr_IF_18 & ((\rfif.rdat2[12]~399_combout  & (\regs[29][12]~q )) # (!\rfif.rdat2[12]~399_combout  & ((\regs[21][12]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[12]~399_combout ))))

	.dataa(\regs[29][12]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[21][12]~q ),
	.datad(\rfif.rdat2[12]~399_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~400_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~400 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[12]~400 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N11
dffeas \regs[28][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][12] .is_wysiwyg = "true";
defparam \regs[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N7
dffeas \regs[16][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][12] .is_wysiwyg = "true";
defparam \regs[16][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N13
dffeas \regs[20][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][12] .is_wysiwyg = "true";
defparam \regs[20][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[12]~403 (
// Equation(s):
// \rfif.rdat2[12]~403_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[20][12]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[16][12]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][12]~q ),
	.datad(\regs[20][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~403_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~403 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[12]~403 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[12]~404 (
// Equation(s):
// \rfif.rdat2[12]~404_combout  = (Instr_IF_19 & ((\rfif.rdat2[12]~403_combout  & ((\regs[28][12]~q ))) # (!\rfif.rdat2[12]~403_combout  & (\regs[24][12]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[12]~403_combout ))))

	.dataa(\regs[24][12]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[28][12]~q ),
	.datad(\rfif.rdat2[12]~403_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~404_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~404 .lut_mask = 16'hF388;
defparam \rfif.rdat2[12]~404 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N9
dffeas \regs[26][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][12] .is_wysiwyg = "true";
defparam \regs[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N11
dffeas \regs[30][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][12] .is_wysiwyg = "true";
defparam \regs[30][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \regs[18][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][12] .is_wysiwyg = "true";
defparam \regs[18][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N29
dffeas \regs[22][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][12] .is_wysiwyg = "true";
defparam \regs[22][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[12]~401 (
// Equation(s):
// \rfif.rdat2[12]~401_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][12]~q ))) # (!Instr_IF_18 & (\regs[18][12]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][12]~q ),
	.datad(\regs[22][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~401_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~401 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[12]~401 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[12]~402 (
// Equation(s):
// \rfif.rdat2[12]~402_combout  = (Instr_IF_19 & ((\rfif.rdat2[12]~401_combout  & ((\regs[30][12]~q ))) # (!\rfif.rdat2[12]~401_combout  & (\regs[26][12]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[12]~401_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][12]~q ),
	.datac(\regs[30][12]~q ),
	.datad(\rfif.rdat2[12]~401_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~402_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~402 .lut_mask = 16'hF588;
defparam \rfif.rdat2[12]~402 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[12]~405 (
// Equation(s):
// \rfif.rdat2[12]~405_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\rfif.rdat2[12]~402_combout )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\rfif.rdat2[12]~404_combout )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[12]~404_combout ),
	.datad(\rfif.rdat2[12]~402_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~405_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~405 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[12]~405 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N5
dffeas \regs[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][12] .is_wysiwyg = "true";
defparam \regs[23][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N31
dffeas \regs[31][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][12] .is_wysiwyg = "true";
defparam \regs[31][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[12]~407 (
// Equation(s):
// \rfif.rdat2[12]~407_combout  = (\rfif.rdat2[12]~406_combout  & (((\regs[31][12]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[12]~406_combout  & (\regs[23][12]~q  & ((Instr_IF_18))))

	.dataa(\rfif.rdat2[12]~406_combout ),
	.datab(\regs[23][12]~q ),
	.datac(\regs[31][12]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~407_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~407 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[12]~407 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[12]~408 (
// Equation(s):
// \rfif.rdat2[12]~408_combout  = (Instr_IF_16 & ((\rfif.rdat2[12]~405_combout  & ((\rfif.rdat2[12]~407_combout ))) # (!\rfif.rdat2[12]~405_combout  & (\rfif.rdat2[12]~400_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[12]~405_combout ))))

	.dataa(\rfif.rdat2[12]~400_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[12]~405_combout ),
	.datad(\rfif.rdat2[12]~407_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~408_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~408 .lut_mask = 16'hF838;
defparam \rfif.rdat2[12]~408 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N31
dffeas \regs[6][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][12] .is_wysiwyg = "true";
defparam \regs[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N1
dffeas \regs[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][12] .is_wysiwyg = "true";
defparam \regs[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \rfif.rdat2[12]~409 (
// Equation(s):
// \rfif.rdat2[12]~409_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[5][12]~q )) # (!Instr_IF_16 & ((\regs[4][12]~q )))))

	.dataa(\regs[5][12]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[4][12]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~409_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~409 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[12]~409 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \rfif.rdat2[12]~410 (
// Equation(s):
// \rfif.rdat2[12]~410_combout  = (Instr_IF_17 & ((\rfif.rdat2[12]~409_combout  & (\regs[7][12]~q )) # (!\rfif.rdat2[12]~409_combout  & ((\regs[6][12]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[12]~409_combout ))))

	.dataa(\regs[7][12]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[6][12]~q ),
	.datad(\rfif.rdat2[12]~409_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~410_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~410 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[12]~410 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N23
dffeas \regs[0][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][12] .is_wysiwyg = "true";
defparam \regs[0][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[12]~413 (
// Equation(s):
// \rfif.rdat2[12]~413_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][12]~q )) # (!Instr_IF_17 & ((\regs[0][12]~q )))))

	.dataa(\regs[2][12]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[0][12]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~413_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~413 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[12]~413 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N5
dffeas \regs[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][12] .is_wysiwyg = "true";
defparam \regs[3][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N7
dffeas \regs[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][12] .is_wysiwyg = "true";
defparam \regs[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \rfif.rdat2[12]~414 (
// Equation(s):
// \rfif.rdat2[12]~414_combout  = (Instr_IF_16 & ((\rfif.rdat2[12]~413_combout  & (\regs[3][12]~q )) # (!\rfif.rdat2[12]~413_combout  & ((\regs[1][12]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[12]~413_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[12]~413_combout ),
	.datac(\regs[3][12]~q ),
	.datad(\regs[1][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~414_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~414 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[12]~414 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N31
dffeas \regs[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][12] .is_wysiwyg = "true";
defparam \regs[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \regs[10][12]~feeder (
// Equation(s):
// \regs[10][12]~feeder_combout  = \input_a~99_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a2),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][12]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N29
dffeas \regs[10][12] (
	.clk(!CLK),
	.d(\regs[10][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][12] .is_wysiwyg = "true";
defparam \regs[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \rfif.rdat2[12]~411 (
// Equation(s):
// \rfif.rdat2[12]~411_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[10][12]~q ))) # (!Instr_IF_17 & (\regs[8][12]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][12]~q ),
	.datad(\regs[10][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~411_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~411 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[12]~411 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N7
dffeas \regs[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][12] .is_wysiwyg = "true";
defparam \regs[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N1
dffeas \regs[9][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][12] .is_wysiwyg = "true";
defparam \regs[9][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \rfif.rdat2[12]~412 (
// Equation(s):
// \rfif.rdat2[12]~412_combout  = (Instr_IF_16 & ((\rfif.rdat2[12]~411_combout  & (\regs[11][12]~q )) # (!\rfif.rdat2[12]~411_combout  & ((\regs[9][12]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[12]~411_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[12]~411_combout ),
	.datac(\regs[11][12]~q ),
	.datad(\regs[9][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~412_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~412 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[12]~412 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[12]~415 (
// Equation(s):
// \rfif.rdat2[12]~415_combout  = (Instr_IF_19 & (((\rfif.rdat2[12]~412_combout ) # (Instr_IF_18)))) # (!Instr_IF_19 & (\rfif.rdat2[12]~414_combout  & ((!Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[12]~414_combout ),
	.datac(\rfif.rdat2[12]~412_combout ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~415_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~415 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[12]~415 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N24
cycloneive_lcell_comb \regs[15][12]~feeder (
// Equation(s):
// \regs[15][12]~feeder_combout  = \input_a~99_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a2),
	.cin(gnd),
	.combout(\regs[15][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y29_N25
dffeas \regs[15][12] (
	.clk(!CLK),
	.d(\regs[15][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][12] .is_wysiwyg = "true";
defparam \regs[15][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \regs[14][12]~feeder (
// Equation(s):
// \regs[14][12]~feeder_combout  = \input_a~99_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a2),
	.cin(gnd),
	.combout(\regs[14][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[14][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N19
dffeas \regs[14][12] (
	.clk(!CLK),
	.d(\regs[14][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][12] .is_wysiwyg = "true";
defparam \regs[14][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[12]~417 (
// Equation(s):
// \rfif.rdat2[12]~417_combout  = (\rfif.rdat2[12]~416_combout  & ((\regs[15][12]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[12]~416_combout  & (((Instr_IF_17 & \regs[14][12]~q ))))

	.dataa(\rfif.rdat2[12]~416_combout ),
	.datab(\regs[15][12]~q ),
	.datac(Instr_IF_17),
	.datad(\regs[14][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~417_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~417 .lut_mask = 16'hDA8A;
defparam \rfif.rdat2[12]~417 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[12]~418 (
// Equation(s):
// \rfif.rdat2[12]~418_combout  = (Instr_IF_18 & ((\rfif.rdat2[12]~415_combout  & ((\rfif.rdat2[12]~417_combout ))) # (!\rfif.rdat2[12]~415_combout  & (\rfif.rdat2[12]~410_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[12]~415_combout ))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[12]~410_combout ),
	.datac(\rfif.rdat2[12]~415_combout ),
	.datad(\rfif.rdat2[12]~417_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[12]~418_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[12]~418 .lut_mask = 16'hF858;
defparam \rfif.rdat2[12]~418 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N25
dffeas \regs[24][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][12] .is_wysiwyg = "true";
defparam \regs[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[12]~384 (
// Equation(s):
// \rfif.rdat1[12]~384_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[24][12]~q )) # (!Instr_IF_24 & ((\regs[16][12]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[24][12]~q ),
	.datad(\regs[16][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~384_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~384 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[12]~384 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[12]~385 (
// Equation(s):
// \rfif.rdat1[12]~385_combout  = (\rfif.rdat1[12]~384_combout  & ((\regs[28][12]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[12]~384_combout  & (((\regs[20][12]~q  & Instr_IF_23))))

	.dataa(\regs[28][12]~q ),
	.datab(\rfif.rdat1[12]~384_combout ),
	.datac(\regs[20][12]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~385_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~385 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[12]~385 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N15
dffeas \regs[29][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][12] .is_wysiwyg = "true";
defparam \regs[29][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N19
dffeas \regs[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][12] .is_wysiwyg = "true";
defparam \regs[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[12]~382 (
// Equation(s):
// \rfif.rdat1[12]~382_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][12]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[17][12]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[17][12]~q ),
	.datad(\regs[21][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~382_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~382 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[12]~382 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[12]~383 (
// Equation(s):
// \rfif.rdat1[12]~383_combout  = (Instr_IF_24 & ((\rfif.rdat1[12]~382_combout  & ((\regs[29][12]~q ))) # (!\rfif.rdat1[12]~382_combout  & (\regs[25][12]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[12]~382_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[25][12]~q ),
	.datac(\regs[29][12]~q ),
	.datad(\rfif.rdat1[12]~382_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~383_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~383 .lut_mask = 16'hF588;
defparam \rfif.rdat1[12]~383 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N24
cycloneive_lcell_comb \rfif.rdat1[12]~386 (
// Equation(s):
// \rfif.rdat1[12]~386_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & ((\rfif.rdat1[12]~383_combout ))) # (!Instr_IF_21 & (\rfif.rdat1[12]~385_combout ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[12]~385_combout ),
	.datad(\rfif.rdat1[12]~383_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~386_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~386 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[12]~386 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[12]~387 (
// Equation(s):
// \rfif.rdat1[12]~387_combout  = (Instr_IF_23 & (((\regs[23][12]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[19][12]~q  & ((!Instr_IF_24))))

	.dataa(\regs[19][12]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[23][12]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~387_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~387 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[12]~387 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N25
dffeas \regs[27][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][12] .is_wysiwyg = "true";
defparam \regs[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[12]~388 (
// Equation(s):
// \rfif.rdat1[12]~388_combout  = (Instr_IF_24 & ((\rfif.rdat1[12]~387_combout  & ((\regs[31][12]~q ))) # (!\rfif.rdat1[12]~387_combout  & (\regs[27][12]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[12]~387_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[12]~387_combout ),
	.datac(\regs[27][12]~q ),
	.datad(\regs[31][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~388_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~388 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[12]~388 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[12]~380 (
// Equation(s):
// \rfif.rdat1[12]~380_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][12]~q )) # (!Instr_IF_24 & ((\regs[18][12]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][12]~q ),
	.datad(\regs[18][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~380_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~380 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[12]~380 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[12]~381 (
// Equation(s):
// \rfif.rdat1[12]~381_combout  = (Instr_IF_23 & ((\rfif.rdat1[12]~380_combout  & (\regs[30][12]~q )) # (!\rfif.rdat1[12]~380_combout  & ((\regs[22][12]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[12]~380_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[30][12]~q ),
	.datac(\regs[22][12]~q ),
	.datad(\rfif.rdat1[12]~380_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~381_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~381 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[12]~381 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[12]~390 (
// Equation(s):
// \rfif.rdat1[12]~390_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[9][12]~q )) # (!Instr_IF_21 & ((\regs[8][12]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[9][12]~q ),
	.datad(\regs[8][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~390_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~390 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[12]~390 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[12]~391 (
// Equation(s):
// \rfif.rdat1[12]~391_combout  = (\rfif.rdat1[12]~390_combout  & ((\regs[11][12]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[12]~390_combout  & (((\regs[10][12]~q  & Instr_IF_22))))

	.dataa(\regs[11][12]~q ),
	.datab(\regs[10][12]~q ),
	.datac(\rfif.rdat1[12]~390_combout ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~391_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~391 .lut_mask = 16'hACF0;
defparam \rfif.rdat1[12]~391 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \regs[2][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][12] .is_wysiwyg = "true";
defparam \regs[2][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[12]~395 (
// Equation(s):
// \rfif.rdat1[12]~395_combout  = (\rfif.rdat1[12]~394_combout  & (((\regs[3][12]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[12]~394_combout  & (Instr_IF_22 & (\regs[2][12]~q )))

	.dataa(\rfif.rdat1[12]~394_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[2][12]~q ),
	.datad(\regs[3][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~395_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~395 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[12]~395 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \regs[5][12]~feeder (
// Equation(s):
// \regs[5][12]~feeder_combout  = \input_a~99_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a2),
	.cin(gnd),
	.combout(\regs[5][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][12]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N29
dffeas \regs[5][12] (
	.clk(!CLK),
	.d(\regs[5][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][12] .is_wysiwyg = "true";
defparam \regs[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \rfif.rdat1[12]~392 (
// Equation(s):
// \rfif.rdat1[12]~392_combout  = (Instr_IF_22 & (((\regs[6][12]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[4][12]~q  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[4][12]~q ),
	.datac(\regs[6][12]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~392_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~392 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[12]~392 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[12]~393 (
// Equation(s):
// \rfif.rdat1[12]~393_combout  = (Instr_IF_21 & ((\rfif.rdat1[12]~392_combout  & (\regs[7][12]~q )) # (!\rfif.rdat1[12]~392_combout  & ((\regs[5][12]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[12]~392_combout ))))

	.dataa(\regs[7][12]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][12]~q ),
	.datad(\rfif.rdat1[12]~392_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~393_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~393 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[12]~393 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[12]~396 (
// Equation(s):
// \rfif.rdat1[12]~396_combout  = (Instr_IF_23 & (((\rfif.rdat1[12]~393_combout ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\rfif.rdat1[12]~395_combout  & ((!Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[12]~395_combout ),
	.datac(\rfif.rdat1[12]~393_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~396_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~396 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[12]~396 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N11
dffeas \regs[12][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][12] .is_wysiwyg = "true";
defparam \regs[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[12]~397 (
// Equation(s):
// \rfif.rdat1[12]~397_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[14][12]~q ))) # (!Instr_IF_22 & (\regs[12][12]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][12]~q ),
	.datac(Instr_IF_22),
	.datad(\regs[14][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~397_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~397 .lut_mask = 16'hF4A4;
defparam \rfif.rdat1[12]~397 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N9
dffeas \regs[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][12] .is_wysiwyg = "true";
defparam \regs[13][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[12]~398 (
// Equation(s):
// \rfif.rdat1[12]~398_combout  = (\rfif.rdat1[12]~397_combout  & (((\regs[15][12]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[12]~397_combout  & (Instr_IF_21 & (\regs[13][12]~q )))

	.dataa(\rfif.rdat1[12]~397_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[13][12]~q ),
	.datad(\regs[15][12]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[12]~398_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[12]~398 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[12]~398 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N20
cycloneive_lcell_comb \regs[11][11]~feeder (
// Equation(s):
// \regs[11][11]~feeder_combout  = \input_a~102_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a3),
	.cin(gnd),
	.combout(\regs[11][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[11][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N21
dffeas \regs[11][11] (
	.clk(!CLK),
	.d(\regs[11][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][11] .is_wysiwyg = "true";
defparam \regs[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N13
dffeas \regs[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][11] .is_wysiwyg = "true";
defparam \regs[10][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N23
dffeas \regs[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][11] .is_wysiwyg = "true";
defparam \regs[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N26
cycloneive_lcell_comb \regs[9][11]~feeder (
// Equation(s):
// \regs[9][11]~feeder_combout  = \input_a~102_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a3),
	.cin(gnd),
	.combout(\regs[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][11]~feeder .lut_mask = 16'hFF00;
defparam \regs[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N27
dffeas \regs[9][11] (
	.clk(!CLK),
	.d(\regs[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][11] .is_wysiwyg = "true";
defparam \regs[9][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[11]~430 (
// Equation(s):
// \rfif.rdat2[11]~430_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][11]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][11]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][11]~q ),
	.datad(\regs[9][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~430_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~430 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[11]~430 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[11]~431 (
// Equation(s):
// \rfif.rdat2[11]~431_combout  = (Instr_IF_17 & ((\rfif.rdat2[11]~430_combout  & (\regs[11][11]~q )) # (!\rfif.rdat2[11]~430_combout  & ((\regs[10][11]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[11]~430_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[11][11]~q ),
	.datac(\regs[10][11]~q ),
	.datad(\rfif.rdat2[11]~430_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~431_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~431 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[11]~431 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N3
dffeas \regs[13][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][11] .is_wysiwyg = "true";
defparam \regs[13][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N1
dffeas \regs[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][11] .is_wysiwyg = "true";
defparam \regs[12][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N13
dffeas \regs[14][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][11] .is_wysiwyg = "true";
defparam \regs[14][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[11]~437 (
// Equation(s):
// \rfif.rdat2[11]~437_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][11]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][11]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][11]~q ),
	.datad(\regs[14][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~437_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~437 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[11]~437 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[11]~438 (
// Equation(s):
// \rfif.rdat2[11]~438_combout  = (Instr_IF_16 & ((\rfif.rdat2[11]~437_combout  & (\regs[15][11]~q )) # (!\rfif.rdat2[11]~437_combout  & ((\regs[13][11]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[11]~437_combout ))))

	.dataa(\regs[15][11]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[13][11]~q ),
	.datad(\rfif.rdat2[11]~437_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~438_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~438 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[11]~438 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N25
dffeas \regs[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][11] .is_wysiwyg = "true";
defparam \regs[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \rfif.rdat2[11]~432 (
// Equation(s):
// \rfif.rdat2[11]~432_combout  = (Instr_IF_17 & ((\regs[6][11]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\regs[4][11]~q  & !Instr_IF_16))))

	.dataa(\regs[6][11]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[4][11]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~432_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~432 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[11]~432 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N31
dffeas \regs[7][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][11] .is_wysiwyg = "true";
defparam \regs[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N13
dffeas \regs[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][11] .is_wysiwyg = "true";
defparam \regs[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[11]~433 (
// Equation(s):
// \rfif.rdat2[11]~433_combout  = (Instr_IF_16 & ((\rfif.rdat2[11]~432_combout  & (\regs[7][11]~q )) # (!\rfif.rdat2[11]~432_combout  & ((\regs[5][11]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[11]~432_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[11]~432_combout ),
	.datac(\regs[7][11]~q ),
	.datad(\regs[5][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~433_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~433 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[11]~433 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[11]~436 (
// Equation(s):
// \rfif.rdat2[11]~436_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & ((\rfif.rdat2[11]~433_combout ))) # (!Instr_IF_18 & (\rfif.rdat2[11]~435_combout ))))

	.dataa(\rfif.rdat2[11]~435_combout ),
	.datab(Instr_IF_19),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[11]~433_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~436_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~436 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[11]~436 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[11]~439 (
// Equation(s):
// \rfif.rdat2[11]~439_combout  = (Instr_IF_19 & ((\rfif.rdat2[11]~436_combout  & ((\rfif.rdat2[11]~438_combout ))) # (!\rfif.rdat2[11]~436_combout  & (\rfif.rdat2[11]~431_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[11]~436_combout ))))

	.dataa(\rfif.rdat2[11]~431_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[11]~438_combout ),
	.datad(\rfif.rdat2[11]~436_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~439_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~439 .lut_mask = 16'hF388;
defparam \rfif.rdat2[11]~439 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N1
dffeas \regs[22][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][11] .is_wysiwyg = "true";
defparam \regs[22][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N15
dffeas \regs[18][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][11] .is_wysiwyg = "true";
defparam \regs[18][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N1
dffeas \regs[26][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][11] .is_wysiwyg = "true";
defparam \regs[26][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \rfif.rdat2[11]~420 (
// Equation(s):
// \rfif.rdat2[11]~420_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[26][11]~q ))) # (!Instr_IF_19 & (\regs[18][11]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[18][11]~q ),
	.datac(\regs[26][11]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~420_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~420 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[11]~420 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \rfif.rdat2[11]~421 (
// Equation(s):
// \rfif.rdat2[11]~421_combout  = (Instr_IF_18 & ((\rfif.rdat2[11]~420_combout  & (\regs[30][11]~q )) # (!\rfif.rdat2[11]~420_combout  & ((\regs[22][11]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[11]~420_combout ))))

	.dataa(\regs[30][11]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][11]~q ),
	.datad(\rfif.rdat2[11]~420_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~421_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~421 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[11]~421 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N1
dffeas \regs[27][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][11] .is_wysiwyg = "true";
defparam \regs[27][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \regs[31][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][11] .is_wysiwyg = "true";
defparam \regs[31][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N21
dffeas \regs[19][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][11] .is_wysiwyg = "true";
defparam \regs[19][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N11
dffeas \regs[23][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][11] .is_wysiwyg = "true";
defparam \regs[23][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[11]~427 (
// Equation(s):
// \rfif.rdat2[11]~427_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[23][11]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[19][11]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][11]~q ),
	.datad(\regs[23][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~427_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~427 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[11]~427 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[11]~428 (
// Equation(s):
// \rfif.rdat2[11]~428_combout  = (Instr_IF_19 & ((\rfif.rdat2[11]~427_combout  & ((\regs[31][11]~q ))) # (!\rfif.rdat2[11]~427_combout  & (\regs[27][11]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[11]~427_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[27][11]~q ),
	.datac(\regs[31][11]~q ),
	.datad(\rfif.rdat2[11]~427_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~428_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~428 .lut_mask = 16'hF588;
defparam \rfif.rdat2[11]~428 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N27
dffeas \regs[28][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][11] .is_wysiwyg = "true";
defparam \regs[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N25
dffeas \regs[20][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][11] .is_wysiwyg = "true";
defparam \regs[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[11]~425 (
// Equation(s):
// \rfif.rdat2[11]~425_combout  = (\rfif.rdat2[11]~424_combout  & (((\regs[28][11]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[11]~424_combout  & (Instr_IF_18 & ((\regs[20][11]~q ))))

	.dataa(\rfif.rdat2[11]~424_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[28][11]~q ),
	.datad(\regs[20][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~425_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~425 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[11]~425 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N5
dffeas \regs[25][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][11] .is_wysiwyg = "true";
defparam \regs[25][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N11
dffeas \regs[29][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][11] .is_wysiwyg = "true";
defparam \regs[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N19
dffeas \regs[17][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][11] .is_wysiwyg = "true";
defparam \regs[17][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N17
dffeas \regs[21][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][11] .is_wysiwyg = "true";
defparam \regs[21][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[11]~422 (
// Equation(s):
// \rfif.rdat2[11]~422_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][11]~q ))) # (!Instr_IF_18 & (\regs[17][11]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][11]~q ),
	.datad(\regs[21][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~422_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~422 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[11]~422 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[11]~423 (
// Equation(s):
// \rfif.rdat2[11]~423_combout  = (Instr_IF_19 & ((\rfif.rdat2[11]~422_combout  & ((\regs[29][11]~q ))) # (!\rfif.rdat2[11]~422_combout  & (\regs[25][11]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[11]~422_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][11]~q ),
	.datac(\regs[29][11]~q ),
	.datad(\rfif.rdat2[11]~422_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~423_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~423 .lut_mask = 16'hF588;
defparam \rfif.rdat2[11]~423 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \rfif.rdat2[11]~426 (
// Equation(s):
// \rfif.rdat2[11]~426_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\rfif.rdat2[11]~423_combout ))) # (!Instr_IF_16 & (\rfif.rdat2[11]~425_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[11]~425_combout ),
	.datac(\rfif.rdat2[11]~423_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~426_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~426 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[11]~426 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[11]~429 (
// Equation(s):
// \rfif.rdat2[11]~429_combout  = (Instr_IF_17 & ((\rfif.rdat2[11]~426_combout  & ((\rfif.rdat2[11]~428_combout ))) # (!\rfif.rdat2[11]~426_combout  & (\rfif.rdat2[11]~421_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[11]~426_combout ))))

	.dataa(\rfif.rdat2[11]~421_combout ),
	.datab(\rfif.rdat2[11]~428_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[11]~426_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[11]~429_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[11]~429 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[11]~429 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[11]~407 (
// Equation(s):
// \rfif.rdat1[11]~407_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[27][11]~q ))) # (!Instr_IF_24 & (\regs[19][11]~q ))))

	.dataa(\regs[19][11]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[27][11]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~407_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~407 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[11]~407 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \rfif.rdat1[11]~408 (
// Equation(s):
// \rfif.rdat1[11]~408_combout  = (Instr_IF_23 & ((\rfif.rdat1[11]~407_combout  & (\regs[31][11]~q )) # (!\rfif.rdat1[11]~407_combout  & ((\regs[23][11]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[11]~407_combout ))))

	.dataa(\regs[31][11]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[23][11]~q ),
	.datad(\rfif.rdat1[11]~407_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~408_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~408 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[11]~408 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[11]~400 (
// Equation(s):
// \rfif.rdat1[11]~400_combout  = (Instr_IF_24 & (((\regs[25][11]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][11]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][11]~q ),
	.datac(\regs[25][11]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~400_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~400 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[11]~400 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[11]~401 (
// Equation(s):
// \rfif.rdat1[11]~401_combout  = (\rfif.rdat1[11]~400_combout  & (((\regs[29][11]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[11]~400_combout  & (Instr_IF_23 & (\regs[21][11]~q )))

	.dataa(\rfif.rdat1[11]~400_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[21][11]~q ),
	.datad(\regs[29][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~401_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~401 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[11]~401 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[11]~404 (
// Equation(s):
// \rfif.rdat1[11]~404_combout  = (Instr_IF_23 & (((\regs[20][11]~q ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\regs[16][11]~q  & ((!Instr_IF_24))))

	.dataa(\regs[16][11]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[20][11]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~404_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~404 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[11]~404 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N25
dffeas \regs[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][11] .is_wysiwyg = "true";
defparam \regs[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[11]~405 (
// Equation(s):
// \rfif.rdat1[11]~405_combout  = (\rfif.rdat1[11]~404_combout  & ((\regs[28][11]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[11]~404_combout  & (((\regs[24][11]~q  & Instr_IF_24))))

	.dataa(\regs[28][11]~q ),
	.datab(\rfif.rdat1[11]~404_combout ),
	.datac(\regs[24][11]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~405_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~405 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[11]~405 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \rfif.rdat1[11]~402 (
// Equation(s):
// \rfif.rdat1[11]~402_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][11]~q ))) # (!Instr_IF_23 & (\regs[18][11]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[18][11]~q ),
	.datad(\regs[22][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~402_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~402 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[11]~402 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N11
dffeas \regs[30][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][11] .is_wysiwyg = "true";
defparam \regs[30][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \rfif.rdat1[11]~403 (
// Equation(s):
// \rfif.rdat1[11]~403_combout  = (Instr_IF_24 & ((\rfif.rdat1[11]~402_combout  & (\regs[30][11]~q )) # (!\rfif.rdat1[11]~402_combout  & ((\regs[26][11]~q ))))) # (!Instr_IF_24 & (\rfif.rdat1[11]~402_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[11]~402_combout ),
	.datac(\regs[30][11]~q ),
	.datad(\regs[26][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~403_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~403 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[11]~403 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \rfif.rdat1[11]~406 (
// Equation(s):
// \rfif.rdat1[11]~406_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[11]~403_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[11]~405_combout ))))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[11]~405_combout ),
	.datac(\rfif.rdat1[11]~403_combout ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~406_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~406 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[11]~406 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \rfif.rdat1[11]~417 (
// Equation(s):
// \rfif.rdat1[11]~417_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[13][11]~q ))) # (!Instr_IF_21 & (\regs[12][11]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[12][11]~q ),
	.datad(\regs[13][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~417_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~417 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[11]~417 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y30_N15
dffeas \regs[15][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][11] .is_wysiwyg = "true";
defparam \regs[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[11]~418 (
// Equation(s):
// \rfif.rdat1[11]~418_combout  = (\rfif.rdat1[11]~417_combout  & (((\regs[15][11]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[11]~417_combout  & (Instr_IF_22 & (\regs[14][11]~q )))

	.dataa(\rfif.rdat1[11]~417_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[14][11]~q ),
	.datad(\regs[15][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~418_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~418 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[11]~418 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[11]~412 (
// Equation(s):
// \rfif.rdat1[11]~412_combout  = (Instr_IF_22 & (((\regs[10][11]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[8][11]~q  & ((!Instr_IF_21))))

	.dataa(\regs[8][11]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[10][11]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~412_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~412 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[11]~412 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N28
cycloneive_lcell_comb \rfif.rdat1[11]~413 (
// Equation(s):
// \rfif.rdat1[11]~413_combout  = (Instr_IF_21 & ((\rfif.rdat1[11]~412_combout  & ((\regs[11][11]~q ))) # (!\rfif.rdat1[11]~412_combout  & (\regs[9][11]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[11]~412_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[11]~412_combout ),
	.datac(\regs[9][11]~q ),
	.datad(\regs[11][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~413_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~413 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[11]~413 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \regs[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][11] .is_wysiwyg = "true";
defparam \regs[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N19
dffeas \regs[0][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][11] .is_wysiwyg = "true";
defparam \regs[0][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[11]~414 (
// Equation(s):
// \rfif.rdat1[11]~414_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[2][11]~q )) # (!Instr_IF_22 & ((\regs[0][11]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[2][11]~q ),
	.datad(\regs[0][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~414_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~414 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[11]~414 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N21
dffeas \regs[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][11] .is_wysiwyg = "true";
defparam \regs[1][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N19
dffeas \regs[3][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][11] .is_wysiwyg = "true";
defparam \regs[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[11]~415 (
// Equation(s):
// \rfif.rdat1[11]~415_combout  = (Instr_IF_21 & ((\rfif.rdat1[11]~414_combout  & ((\regs[3][11]~q ))) # (!\rfif.rdat1[11]~414_combout  & (\regs[1][11]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[11]~414_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[11]~414_combout ),
	.datac(\regs[1][11]~q ),
	.datad(\regs[3][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~415_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~415 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[11]~415 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[11]~416 (
// Equation(s):
// \rfif.rdat1[11]~416_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & (\rfif.rdat1[11]~413_combout )) # (!Instr_IF_24 & ((\rfif.rdat1[11]~415_combout )))))

	.dataa(\rfif.rdat1[11]~413_combout ),
	.datab(Instr_IF_23),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[11]~415_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~416_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~416 .lut_mask = 16'hE3E0;
defparam \rfif.rdat1[11]~416 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N11
dffeas \regs[6][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][11] .is_wysiwyg = "true";
defparam \regs[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[11]~410 (
// Equation(s):
// \rfif.rdat1[11]~410_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[5][11]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[4][11]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[5][11]~q ),
	.datad(\regs[4][11]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~410_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~410 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[11]~410 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \rfif.rdat1[11]~411 (
// Equation(s):
// \rfif.rdat1[11]~411_combout  = (Instr_IF_22 & ((\rfif.rdat1[11]~410_combout  & (\regs[7][11]~q )) # (!\rfif.rdat1[11]~410_combout  & ((\regs[6][11]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[11]~410_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[7][11]~q ),
	.datac(\regs[6][11]~q ),
	.datad(\rfif.rdat1[11]~410_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[11]~411_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[11]~411 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[11]~411 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N5
dffeas \regs[13][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][10] .is_wysiwyg = "true";
defparam \regs[13][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N7
dffeas \regs[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][10] .is_wysiwyg = "true";
defparam \regs[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \rfif.rdat2[10]~458 (
// Equation(s):
// \rfif.rdat2[10]~458_combout  = (Instr_IF_16 & ((\regs[13][10]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[12][10]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[13][10]~q ),
	.datac(\regs[12][10]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~458_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~458 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[10]~458 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N21
dffeas \regs[14][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][10] .is_wysiwyg = "true";
defparam \regs[14][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \regs[15][10]~feeder (
// Equation(s):
// \regs[15][10]~feeder_combout  = \input_a~105_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a4),
	.cin(gnd),
	.combout(\regs[15][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][10]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N17
dffeas \regs[15][10] (
	.clk(!CLK),
	.d(\regs[15][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][10] .is_wysiwyg = "true";
defparam \regs[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[10]~459 (
// Equation(s):
// \rfif.rdat2[10]~459_combout  = (Instr_IF_17 & ((\rfif.rdat2[10]~458_combout  & ((\regs[15][10]~q ))) # (!\rfif.rdat2[10]~458_combout  & (\regs[14][10]~q )))) # (!Instr_IF_17 & (\rfif.rdat2[10]~458_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[10]~458_combout ),
	.datac(\regs[14][10]~q ),
	.datad(\regs[15][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~459_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~459 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[10]~459 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N27
dffeas \regs[6][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][10] .is_wysiwyg = "true";
defparam \regs[6][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N1
dffeas \regs[7][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][10] .is_wysiwyg = "true";
defparam \regs[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N25
dffeas \regs[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][10] .is_wysiwyg = "true";
defparam \regs[4][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N7
dffeas \regs[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][10] .is_wysiwyg = "true";
defparam \regs[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \rfif.rdat2[10]~451 (
// Equation(s):
// \rfif.rdat2[10]~451_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][10]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][10]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][10]~q ),
	.datad(\regs[5][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~451_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~451 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[10]~451 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \rfif.rdat2[10]~452 (
// Equation(s):
// \rfif.rdat2[10]~452_combout  = (Instr_IF_17 & ((\rfif.rdat2[10]~451_combout  & ((\regs[7][10]~q ))) # (!\rfif.rdat2[10]~451_combout  & (\regs[6][10]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[10]~451_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[6][10]~q ),
	.datac(\regs[7][10]~q ),
	.datad(\rfif.rdat2[10]~451_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~452_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~452 .lut_mask = 16'hF588;
defparam \rfif.rdat2[10]~452 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N25
dffeas \regs[9][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][10] .is_wysiwyg = "true";
defparam \regs[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N19
dffeas \regs[11][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][10] .is_wysiwyg = "true";
defparam \regs[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N19
dffeas \regs[8][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][10] .is_wysiwyg = "true";
defparam \regs[8][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N25
dffeas \regs[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][10] .is_wysiwyg = "true";
defparam \regs[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \rfif.rdat2[10]~453 (
// Equation(s):
// \rfif.rdat2[10]~453_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[10][10]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[8][10]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[8][10]~q ),
	.datad(\regs[10][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~453_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~453 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[10]~453 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \rfif.rdat2[10]~454 (
// Equation(s):
// \rfif.rdat2[10]~454_combout  = (Instr_IF_16 & ((\rfif.rdat2[10]~453_combout  & ((\regs[11][10]~q ))) # (!\rfif.rdat2[10]~453_combout  & (\regs[9][10]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[10]~453_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][10]~q ),
	.datac(\regs[11][10]~q ),
	.datad(\rfif.rdat2[10]~453_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~454_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~454 .lut_mask = 16'hF588;
defparam \rfif.rdat2[10]~454 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \rfif.rdat2[10]~457 (
// Equation(s):
// \rfif.rdat2[10]~457_combout  = (Instr_IF_19 & (((Instr_IF_18) # (\rfif.rdat2[10]~454_combout )))) # (!Instr_IF_19 & (\rfif.rdat2[10]~456_combout  & (!Instr_IF_18)))

	.dataa(\rfif.rdat2[10]~456_combout ),
	.datab(Instr_IF_19),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[10]~454_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~457_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~457 .lut_mask = 16'hCEC2;
defparam \rfif.rdat2[10]~457 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[10]~460 (
// Equation(s):
// \rfif.rdat2[10]~460_combout  = (Instr_IF_18 & ((\rfif.rdat2[10]~457_combout  & (\rfif.rdat2[10]~459_combout )) # (!\rfif.rdat2[10]~457_combout  & ((\rfif.rdat2[10]~452_combout ))))) # (!Instr_IF_18 & (((\rfif.rdat2[10]~457_combout ))))

	.dataa(\rfif.rdat2[10]~459_combout ),
	.datab(\rfif.rdat2[10]~452_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[10]~457_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~460_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~460 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[10]~460 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \regs[25][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][10] .is_wysiwyg = "true";
defparam \regs[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N3
dffeas \regs[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][10] .is_wysiwyg = "true";
defparam \regs[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \rfif.rdat2[10]~441 (
// Equation(s):
// \rfif.rdat2[10]~441_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[25][10]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\regs[17][10]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[25][10]~q ),
	.datad(\regs[17][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~441_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~441 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[10]~441 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N1
dffeas \regs[21][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][10] .is_wysiwyg = "true";
defparam \regs[21][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N17
dffeas \regs[29][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][10] .is_wysiwyg = "true";
defparam \regs[29][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \rfif.rdat2[10]~442 (
// Equation(s):
// \rfif.rdat2[10]~442_combout  = (Instr_IF_18 & ((\rfif.rdat2[10]~441_combout  & ((\regs[29][10]~q ))) # (!\rfif.rdat2[10]~441_combout  & (\regs[21][10]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[10]~441_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[10]~441_combout ),
	.datac(\regs[21][10]~q ),
	.datad(\regs[29][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~442_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~442 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[10]~442 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N29
dffeas \regs[19][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][10] .is_wysiwyg = "true";
defparam \regs[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \regs[27][10]~feeder (
// Equation(s):
// \regs[27][10]~feeder_combout  = \input_a~105_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a4),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][10]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N15
dffeas \regs[27][10] (
	.clk(!CLK),
	.d(\regs[27][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][10] .is_wysiwyg = "true";
defparam \regs[27][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[10]~448 (
// Equation(s):
// \rfif.rdat2[10]~448_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[27][10]~q ))) # (!Instr_IF_19 & (\regs[19][10]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][10]~q ),
	.datad(\regs[27][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~448_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~448 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[10]~448 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N31
dffeas \regs[23][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][10] .is_wysiwyg = "true";
defparam \regs[23][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[10]~449 (
// Equation(s):
// \rfif.rdat2[10]~449_combout  = (\rfif.rdat2[10]~448_combout  & ((\regs[31][10]~q ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[10]~448_combout  & (((\regs[23][10]~q  & Instr_IF_18))))

	.dataa(\regs[31][10]~q ),
	.datab(\rfif.rdat2[10]~448_combout ),
	.datac(\regs[23][10]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~449_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~449 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[10]~449 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N31
dffeas \regs[28][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][10] .is_wysiwyg = "true";
defparam \regs[28][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N15
dffeas \regs[16][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][10] .is_wysiwyg = "true";
defparam \regs[16][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N9
dffeas \regs[20][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][10] .is_wysiwyg = "true";
defparam \regs[20][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[10]~445 (
// Equation(s):
// \rfif.rdat2[10]~445_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[20][10]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[16][10]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][10]~q ),
	.datad(\regs[20][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~445_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~445 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[10]~445 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[10]~446 (
// Equation(s):
// \rfif.rdat2[10]~446_combout  = (Instr_IF_19 & ((\rfif.rdat2[10]~445_combout  & ((\regs[28][10]~q ))) # (!\rfif.rdat2[10]~445_combout  & (\regs[24][10]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[10]~445_combout ))))

	.dataa(\regs[24][10]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[28][10]~q ),
	.datad(\rfif.rdat2[10]~445_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~446_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~446 .lut_mask = 16'hF388;
defparam \rfif.rdat2[10]~446 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N15
dffeas \regs[18][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][10] .is_wysiwyg = "true";
defparam \regs[18][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N1
dffeas \regs[22][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][10] .is_wysiwyg = "true";
defparam \regs[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[10]~443 (
// Equation(s):
// \rfif.rdat2[10]~443_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][10]~q ))) # (!Instr_IF_18 & (\regs[18][10]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][10]~q ),
	.datad(\regs[22][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~443_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~443 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[10]~443 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N23
dffeas \regs[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][10] .is_wysiwyg = "true";
defparam \regs[30][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N17
dffeas \regs[26][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][10] .is_wysiwyg = "true";
defparam \regs[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[10]~444 (
// Equation(s):
// \rfif.rdat2[10]~444_combout  = (Instr_IF_19 & ((\rfif.rdat2[10]~443_combout  & (\regs[30][10]~q )) # (!\rfif.rdat2[10]~443_combout  & ((\regs[26][10]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[10]~443_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[10]~443_combout ),
	.datac(\regs[30][10]~q ),
	.datad(\regs[26][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~444_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~444 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[10]~444 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \rfif.rdat2[10]~447 (
// Equation(s):
// \rfif.rdat2[10]~447_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\rfif.rdat2[10]~444_combout )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\rfif.rdat2[10]~446_combout )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[10]~446_combout ),
	.datad(\rfif.rdat2[10]~444_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~447_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~447 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[10]~447 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[10]~450 (
// Equation(s):
// \rfif.rdat2[10]~450_combout  = (Instr_IF_16 & ((\rfif.rdat2[10]~447_combout  & ((\rfif.rdat2[10]~449_combout ))) # (!\rfif.rdat2[10]~447_combout  & (\rfif.rdat2[10]~442_combout )))) # (!Instr_IF_16 & (((\rfif.rdat2[10]~447_combout ))))

	.dataa(\rfif.rdat2[10]~442_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[10]~449_combout ),
	.datad(\rfif.rdat2[10]~447_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[10]~450_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[10]~450 .lut_mask = 16'hF388;
defparam \rfif.rdat2[10]~450 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \rfif.rdat1[10]~427 (
// Equation(s):
// \rfif.rdat1[10]~427_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][10]~q ))) # (!Instr_IF_23 & (\regs[19][10]~q ))))

	.dataa(Instr_IF_24),
	.datab(\regs[19][10]~q ),
	.datac(\regs[23][10]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~427_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~427 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[10]~427 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \regs[31][10]~feeder (
// Equation(s):
// \regs[31][10]~feeder_combout  = \input_a~105_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a4),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[31][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][10]~feeder .lut_mask = 16'hF0F0;
defparam \regs[31][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N27
dffeas \regs[31][10] (
	.clk(!CLK),
	.d(\regs[31][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][10] .is_wysiwyg = "true";
defparam \regs[31][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \rfif.rdat1[10]~428 (
// Equation(s):
// \rfif.rdat1[10]~428_combout  = (\rfif.rdat1[10]~427_combout  & (((\regs[31][10]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[10]~427_combout  & (Instr_IF_24 & (\regs[27][10]~q )))

	.dataa(\rfif.rdat1[10]~427_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[27][10]~q ),
	.datad(\regs[31][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~428_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~428 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[10]~428 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[10]~420 (
// Equation(s):
// \rfif.rdat1[10]~420_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[26][10]~q ))) # (!Instr_IF_24 & (\regs[18][10]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[18][10]~q ),
	.datac(\regs[26][10]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~420_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~420 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[10]~420 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[10]~421 (
// Equation(s):
// \rfif.rdat1[10]~421_combout  = (\rfif.rdat1[10]~420_combout  & ((\regs[30][10]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[10]~420_combout  & (((\regs[22][10]~q  & Instr_IF_23))))

	.dataa(\rfif.rdat1[10]~420_combout ),
	.datab(\regs[30][10]~q ),
	.datac(\regs[22][10]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~421_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~421 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[10]~421 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N1
dffeas \regs[24][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][10] .is_wysiwyg = "true";
defparam \regs[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[10]~424 (
// Equation(s):
// \rfif.rdat1[10]~424_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][10]~q ))) # (!Instr_IF_24 & (\regs[16][10]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][10]~q ),
	.datac(\regs[24][10]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~424_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~424 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[10]~424 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[10]~425 (
// Equation(s):
// \rfif.rdat1[10]~425_combout  = (\rfif.rdat1[10]~424_combout  & ((\regs[28][10]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[10]~424_combout  & (((\regs[20][10]~q  & Instr_IF_23))))

	.dataa(\regs[28][10]~q ),
	.datab(\rfif.rdat1[10]~424_combout ),
	.datac(\regs[20][10]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~425_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~425 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[10]~425 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[10]~422 (
// Equation(s):
// \rfif.rdat1[10]~422_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][10]~q ))) # (!Instr_IF_23 & (\regs[17][10]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[17][10]~q ),
	.datad(\regs[21][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~422_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~422 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[10]~422 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \rfif.rdat1[10]~423 (
// Equation(s):
// \rfif.rdat1[10]~423_combout  = (Instr_IF_24 & ((\rfif.rdat1[10]~422_combout  & (\regs[29][10]~q )) # (!\rfif.rdat1[10]~422_combout  & ((\regs[25][10]~q ))))) # (!Instr_IF_24 & (\rfif.rdat1[10]~422_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[10]~422_combout ),
	.datac(\regs[29][10]~q ),
	.datad(\regs[25][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~423_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~423 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[10]~423 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \rfif.rdat1[10]~426 (
// Equation(s):
// \rfif.rdat1[10]~426_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\rfif.rdat1[10]~423_combout ))) # (!Instr_IF_21 & (\rfif.rdat1[10]~425_combout ))))

	.dataa(\rfif.rdat1[10]~425_combout ),
	.datab(\rfif.rdat1[10]~423_combout ),
	.datac(Instr_IF_22),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~426_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~426 .lut_mask = 16'hFC0A;
defparam \rfif.rdat1[10]~426 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \rfif.rdat1[10]~437 (
// Equation(s):
// \rfif.rdat1[10]~437_combout  = (Instr_IF_22 & ((\regs[14][10]~q ) # ((Instr_IF_21)))) # (!Instr_IF_22 & (((\regs[12][10]~q  & !Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[14][10]~q ),
	.datac(\regs[12][10]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~437_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~437 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[10]~437 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[10]~438 (
// Equation(s):
// \rfif.rdat1[10]~438_combout  = (\rfif.rdat1[10]~437_combout  & (((\regs[15][10]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[10]~437_combout  & (Instr_IF_21 & (\regs[13][10]~q )))

	.dataa(\rfif.rdat1[10]~437_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[13][10]~q ),
	.datad(\regs[15][10]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~438_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~438 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[10]~438 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \rfif.rdat1[10]~433 (
// Equation(s):
// \rfif.rdat1[10]~433_combout  = (\rfif.rdat1[10]~432_combout  & ((\regs[7][10]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[10]~432_combout  & (((\regs[5][10]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[10]~432_combout ),
	.datab(\regs[7][10]~q ),
	.datac(\regs[5][10]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~433_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~433 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[10]~433 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N27
dffeas \regs[3][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][10] .is_wysiwyg = "true";
defparam \regs[3][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N25
dffeas \regs[2][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][10] .is_wysiwyg = "true";
defparam \regs[2][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[10]~435 (
// Equation(s):
// \rfif.rdat1[10]~435_combout  = (\rfif.rdat1[10]~434_combout  & ((\regs[3][10]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[10]~434_combout  & (((\regs[2][10]~q  & Instr_IF_22))))

	.dataa(\rfif.rdat1[10]~434_combout ),
	.datab(\regs[3][10]~q ),
	.datac(\regs[2][10]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~435_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~435 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[10]~435 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N2
cycloneive_lcell_comb \rfif.rdat1[10]~436 (
// Equation(s):
// \rfif.rdat1[10]~436_combout  = (Instr_IF_23 & ((\rfif.rdat1[10]~433_combout ) # ((Instr_IF_24)))) # (!Instr_IF_23 & (((\rfif.rdat1[10]~435_combout  & !Instr_IF_24))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[10]~433_combout ),
	.datac(\rfif.rdat1[10]~435_combout ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~436_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~436 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[10]~436 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[10]~430 (
// Equation(s):
// \rfif.rdat1[10]~430_combout  = (Instr_IF_21 & (((\regs[9][10]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[8][10]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[8][10]~q ),
	.datac(\regs[9][10]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~430_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~430 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[10]~430 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[10]~431 (
// Equation(s):
// \rfif.rdat1[10]~431_combout  = (Instr_IF_22 & ((\rfif.rdat1[10]~430_combout  & (\regs[11][10]~q )) # (!\rfif.rdat1[10]~430_combout  & ((\regs[10][10]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[10]~430_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[11][10]~q ),
	.datac(\regs[10][10]~q ),
	.datad(\rfif.rdat1[10]~430_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[10]~431_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[10]~431 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[10]~431 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N21
dffeas \regs[25][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][9] .is_wysiwyg = "true";
defparam \regs[25][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N7
dffeas \regs[29][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][9] .is_wysiwyg = "true";
defparam \regs[29][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[9]~465 (
// Equation(s):
// \rfif.rdat2[9]~465_combout  = (\rfif.rdat2[9]~464_combout  & (((\regs[29][9]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[9]~464_combout  & (\regs[25][9]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[9]~464_combout ),
	.datab(\regs[25][9]~q ),
	.datac(\regs[29][9]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~465_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~465 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[9]~465 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N11
dffeas \regs[28][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][9] .is_wysiwyg = "true";
defparam \regs[28][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N23
dffeas \regs[16][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][9] .is_wysiwyg = "true";
defparam \regs[16][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N1
dffeas \regs[24][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][9] .is_wysiwyg = "true";
defparam \regs[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[9]~466 (
// Equation(s):
// \rfif.rdat2[9]~466_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][9]~q ))) # (!Instr_IF_19 & (\regs[16][9]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][9]~q ),
	.datad(\regs[24][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~466_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~466 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[9]~466 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[9]~467 (
// Equation(s):
// \rfif.rdat2[9]~467_combout  = (Instr_IF_18 & ((\rfif.rdat2[9]~466_combout  & ((\regs[28][9]~q ))) # (!\rfif.rdat2[9]~466_combout  & (\regs[20][9]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[9]~466_combout ))))

	.dataa(\regs[20][9]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][9]~q ),
	.datad(\rfif.rdat2[9]~466_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~467_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~467 .lut_mask = 16'hF388;
defparam \rfif.rdat2[9]~467 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[9]~468 (
// Equation(s):
// \rfif.rdat2[9]~468_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[9]~465_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[9]~467_combout )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[9]~465_combout ),
	.datad(\rfif.rdat2[9]~467_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~468_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~468 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[9]~468 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N25
dffeas \regs[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][9] .is_wysiwyg = "true";
defparam \regs[22][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N7
dffeas \regs[30][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][9] .is_wysiwyg = "true";
defparam \regs[30][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \rfif.rdat2[9]~463 (
// Equation(s):
// \rfif.rdat2[9]~463_combout  = (\rfif.rdat2[9]~462_combout  & (((\regs[30][9]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[9]~462_combout  & (Instr_IF_18 & (\regs[22][9]~q )))

	.dataa(\rfif.rdat2[9]~462_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[22][9]~q ),
	.datad(\regs[30][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~463_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~463 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[9]~463 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N15
dffeas \regs[31][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][9] .is_wysiwyg = "true";
defparam \regs[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N15
dffeas \regs[23][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][9] .is_wysiwyg = "true";
defparam \regs[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas \regs[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][9] .is_wysiwyg = "true";
defparam \regs[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[9]~469 (
// Equation(s):
// \rfif.rdat2[9]~469_combout  = (Instr_IF_18 & ((\regs[23][9]~q ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((\regs[19][9]~q  & !Instr_IF_19))))

	.dataa(Instr_IF_18),
	.datab(\regs[23][9]~q ),
	.datac(\regs[19][9]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~469_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~469 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[9]~469 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[9]~470 (
// Equation(s):
// \rfif.rdat2[9]~470_combout  = (Instr_IF_19 & ((\rfif.rdat2[9]~469_combout  & ((\regs[31][9]~q ))) # (!\rfif.rdat2[9]~469_combout  & (\regs[27][9]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[9]~469_combout ))))

	.dataa(\regs[27][9]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[31][9]~q ),
	.datad(\rfif.rdat2[9]~469_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~470_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~470 .lut_mask = 16'hF388;
defparam \rfif.rdat2[9]~470 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[9]~471 (
// Equation(s):
// \rfif.rdat2[9]~471_combout  = (Instr_IF_17 & ((\rfif.rdat2[9]~468_combout  & ((\rfif.rdat2[9]~470_combout ))) # (!\rfif.rdat2[9]~468_combout  & (\rfif.rdat2[9]~463_combout )))) # (!Instr_IF_17 & (\rfif.rdat2[9]~468_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[9]~468_combout ),
	.datac(\rfif.rdat2[9]~463_combout ),
	.datad(\rfif.rdat2[9]~470_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~471_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~471 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[9]~471 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N0
cycloneive_lcell_comb \regs[11][9]~feeder (
// Equation(s):
// \regs[11][9]~feeder_combout  = \input_a~108_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a5),
	.cin(gnd),
	.combout(\regs[11][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][9]~feeder .lut_mask = 16'hFF00;
defparam \regs[11][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N1
dffeas \regs[11][9] (
	.clk(!CLK),
	.d(\regs[11][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][9] .is_wysiwyg = "true";
defparam \regs[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N1
dffeas \regs[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][9] .is_wysiwyg = "true";
defparam \regs[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[9]~473 (
// Equation(s):
// \rfif.rdat2[9]~473_combout  = (\rfif.rdat2[9]~472_combout  & ((\regs[11][9]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[9]~472_combout  & (((\regs[10][9]~q  & Instr_IF_17))))

	.dataa(\rfif.rdat2[9]~472_combout ),
	.datab(\regs[11][9]~q ),
	.datac(\regs[10][9]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~473_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~473 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[9]~473 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N19
dffeas \regs[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][9] .is_wysiwyg = "true";
defparam \regs[13][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N17
dffeas \regs[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][9] .is_wysiwyg = "true";
defparam \regs[12][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N1
dffeas \regs[14][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][9] .is_wysiwyg = "true";
defparam \regs[14][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[9]~479 (
// Equation(s):
// \rfif.rdat2[9]~479_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][9]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][9]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][9]~q ),
	.datad(\regs[14][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~479_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~479 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[9]~479 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \rfif.rdat2[9]~480 (
// Equation(s):
// \rfif.rdat2[9]~480_combout  = (Instr_IF_16 & ((\rfif.rdat2[9]~479_combout  & (\regs[15][9]~q )) # (!\rfif.rdat2[9]~479_combout  & ((\regs[13][9]~q ))))) # (!Instr_IF_16 & (((\rfif.rdat2[9]~479_combout ))))

	.dataa(\regs[15][9]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[13][9]~q ),
	.datad(\rfif.rdat2[9]~479_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~480_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~480 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[9]~480 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N9
dffeas \regs[2][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][9] .is_wysiwyg = "true";
defparam \regs[2][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N3
dffeas \regs[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][9] .is_wysiwyg = "true";
defparam \regs[3][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N3
dffeas \regs[0][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][9] .is_wysiwyg = "true";
defparam \regs[0][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \rfif.rdat2[9]~476 (
// Equation(s):
// \rfif.rdat2[9]~476_combout  = (Instr_IF_16 & ((\regs[1][9]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[0][9]~q  & !Instr_IF_17))))

	.dataa(\regs[1][9]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[0][9]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~476_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~476 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[9]~476 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \rfif.rdat2[9]~477 (
// Equation(s):
// \rfif.rdat2[9]~477_combout  = (Instr_IF_17 & ((\rfif.rdat2[9]~476_combout  & ((\regs[3][9]~q ))) # (!\rfif.rdat2[9]~476_combout  & (\regs[2][9]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[9]~476_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[2][9]~q ),
	.datac(\regs[3][9]~q ),
	.datad(\rfif.rdat2[9]~476_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~477_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~477 .lut_mask = 16'hF588;
defparam \rfif.rdat2[9]~477 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N5
dffeas \regs[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][9] .is_wysiwyg = "true";
defparam \regs[5][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N15
dffeas \regs[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][9] .is_wysiwyg = "true";
defparam \regs[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N7
dffeas \regs[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][9] .is_wysiwyg = "true";
defparam \regs[4][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N29
dffeas \regs[6][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][9] .is_wysiwyg = "true";
defparam \regs[6][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[9]~474 (
// Equation(s):
// \rfif.rdat2[9]~474_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][9]~q ))) # (!Instr_IF_17 & (\regs[4][9]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][9]~q ),
	.datad(\regs[6][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~474_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~474 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[9]~474 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[9]~475 (
// Equation(s):
// \rfif.rdat2[9]~475_combout  = (Instr_IF_16 & ((\rfif.rdat2[9]~474_combout  & ((\regs[7][9]~q ))) # (!\rfif.rdat2[9]~474_combout  & (\regs[5][9]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[9]~474_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][9]~q ),
	.datac(\regs[7][9]~q ),
	.datad(\rfif.rdat2[9]~474_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~475_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~475 .lut_mask = 16'hF588;
defparam \rfif.rdat2[9]~475 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[9]~478 (
// Equation(s):
// \rfif.rdat2[9]~478_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\rfif.rdat2[9]~475_combout ))) # (!Instr_IF_18 & (\rfif.rdat2[9]~477_combout ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[9]~477_combout ),
	.datad(\rfif.rdat2[9]~475_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~478_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~478 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[9]~478 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[9]~481 (
// Equation(s):
// \rfif.rdat2[9]~481_combout  = (\rfif.rdat2[9]~478_combout  & (((\rfif.rdat2[9]~480_combout ) # (!Instr_IF_19)))) # (!\rfif.rdat2[9]~478_combout  & (\rfif.rdat2[9]~473_combout  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[9]~473_combout ),
	.datab(\rfif.rdat2[9]~480_combout ),
	.datac(\rfif.rdat2[9]~478_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[9]~481_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[9]~481 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[9]~481 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N1
dffeas \regs[21][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][9] .is_wysiwyg = "true";
defparam \regs[21][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N31
dffeas \regs[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][9] .is_wysiwyg = "true";
defparam \regs[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \rfif.rdat1[9]~440 (
// Equation(s):
// \rfif.rdat1[9]~440_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][9]~q ))) # (!Instr_IF_24 & (\regs[17][9]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[17][9]~q ),
	.datac(\regs[25][9]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~440_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~440 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[9]~440 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \rfif.rdat1[9]~441 (
// Equation(s):
// \rfif.rdat1[9]~441_combout  = (Instr_IF_23 & ((\rfif.rdat1[9]~440_combout  & (\regs[29][9]~q )) # (!\rfif.rdat1[9]~440_combout  & ((\regs[21][9]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[9]~440_combout ))))

	.dataa(\regs[29][9]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[21][9]~q ),
	.datad(\rfif.rdat1[9]~440_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~441_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~441 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[9]~441 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas \regs[27][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][9] .is_wysiwyg = "true";
defparam \regs[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[9]~447 (
// Equation(s):
// \rfif.rdat1[9]~447_combout  = (Instr_IF_24 & (((\regs[27][9]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[19][9]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[19][9]~q ),
	.datac(\regs[27][9]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~447_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~447 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[9]~447 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \rfif.rdat1[9]~448 (
// Equation(s):
// \rfif.rdat1[9]~448_combout  = (\rfif.rdat1[9]~447_combout  & ((\regs[31][9]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[9]~447_combout  & (((\regs[23][9]~q  & Instr_IF_23))))

	.dataa(\regs[31][9]~q ),
	.datab(\rfif.rdat1[9]~447_combout ),
	.datac(\regs[23][9]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~448_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~448 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[9]~448 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[9]~445 (
// Equation(s):
// \rfif.rdat1[9]~445_combout  = (\rfif.rdat1[9]~444_combout  & (((\regs[28][9]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[9]~444_combout  & (Instr_IF_24 & (\regs[24][9]~q )))

	.dataa(\rfif.rdat1[9]~444_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[24][9]~q ),
	.datad(\regs[28][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~445_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~445 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[9]~445 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N5
dffeas \regs[26][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][9] .is_wysiwyg = "true";
defparam \regs[26][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N3
dffeas \regs[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][9] .is_wysiwyg = "true";
defparam \regs[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \rfif.rdat1[9]~442 (
// Equation(s):
// \rfif.rdat1[9]~442_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][9]~q ))) # (!Instr_IF_23 & (\regs[18][9]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[18][9]~q ),
	.datad(\regs[22][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~442_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~442 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[9]~442 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \rfif.rdat1[9]~443 (
// Equation(s):
// \rfif.rdat1[9]~443_combout  = (Instr_IF_24 & ((\rfif.rdat1[9]~442_combout  & ((\regs[30][9]~q ))) # (!\rfif.rdat1[9]~442_combout  & (\regs[26][9]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[9]~442_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[26][9]~q ),
	.datac(\regs[30][9]~q ),
	.datad(\rfif.rdat1[9]~442_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~443_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~443 .lut_mask = 16'hF588;
defparam \rfif.rdat1[9]~443 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[9]~446 (
// Equation(s):
// \rfif.rdat1[9]~446_combout  = (Instr_IF_22 & (((\rfif.rdat1[9]~443_combout ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\rfif.rdat1[9]~445_combout  & ((!Instr_IF_21))))

	.dataa(\rfif.rdat1[9]~445_combout ),
	.datab(\rfif.rdat1[9]~443_combout ),
	.datac(Instr_IF_22),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~446_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~446 .lut_mask = 16'hF0CA;
defparam \rfif.rdat1[9]~446 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N13
dffeas \regs[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][9] .is_wysiwyg = "true";
defparam \regs[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[9]~455 (
// Equation(s):
// \rfif.rdat1[9]~455_combout  = (\rfif.rdat1[9]~454_combout  & ((\regs[3][9]~q ) # ((!Instr_IF_21)))) # (!\rfif.rdat1[9]~454_combout  & (((\regs[1][9]~q  & Instr_IF_21))))

	.dataa(\rfif.rdat1[9]~454_combout ),
	.datab(\regs[3][9]~q ),
	.datac(\regs[1][9]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~455_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~455 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[9]~455 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N0
cycloneive_lcell_comb \rfif.rdat1[9]~452 (
// Equation(s):
// \rfif.rdat1[9]~452_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[10][9]~q ))) # (!Instr_IF_22 & (\regs[8][9]~q ))))

	.dataa(\regs[8][9]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[10][9]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~452_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~452 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[9]~452 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[9]~453 (
// Equation(s):
// \rfif.rdat1[9]~453_combout  = (Instr_IF_21 & ((\rfif.rdat1[9]~452_combout  & ((\regs[11][9]~q ))) # (!\rfif.rdat1[9]~452_combout  & (\regs[9][9]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[9]~452_combout ))))

	.dataa(\regs[9][9]~q ),
	.datab(\regs[11][9]~q ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[9]~452_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~453_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~453 .lut_mask = 16'hCFA0;
defparam \rfif.rdat1[9]~453 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[9]~456 (
// Equation(s):
// \rfif.rdat1[9]~456_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[9]~453_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[9]~455_combout ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[9]~455_combout ),
	.datad(\rfif.rdat1[9]~453_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~456_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~456 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[9]~456 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N29
dffeas \regs[15][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][9] .is_wysiwyg = "true";
defparam \regs[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \rfif.rdat1[9]~457 (
// Equation(s):
// \rfif.rdat1[9]~457_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[13][9]~q )) # (!Instr_IF_21 & ((\regs[12][9]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[13][9]~q ),
	.datad(\regs[12][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~457_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~457 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[9]~457 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[9]~458 (
// Equation(s):
// \rfif.rdat1[9]~458_combout  = (Instr_IF_22 & ((\rfif.rdat1[9]~457_combout  & (\regs[15][9]~q )) # (!\rfif.rdat1[9]~457_combout  & ((\regs[14][9]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[9]~457_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[15][9]~q ),
	.datac(\regs[14][9]~q ),
	.datad(\rfif.rdat1[9]~457_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~458_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~458 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[9]~458 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[9]~450 (
// Equation(s):
// \rfif.rdat1[9]~450_combout  = (Instr_IF_21 & (((\regs[5][9]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[4][9]~q  & ((!Instr_IF_22))))

	.dataa(\regs[4][9]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][9]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~450_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~450 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[9]~450 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[9]~451 (
// Equation(s):
// \rfif.rdat1[9]~451_combout  = (Instr_IF_22 & ((\rfif.rdat1[9]~450_combout  & ((\regs[7][9]~q ))) # (!\rfif.rdat1[9]~450_combout  & (\regs[6][9]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[9]~450_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[9]~450_combout ),
	.datac(\regs[6][9]~q ),
	.datad(\regs[7][9]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[9]~451_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[9]~451 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[9]~451 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N19
dffeas \regs[25][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][8] .is_wysiwyg = "true";
defparam \regs[25][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N15
dffeas \regs[17][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][8] .is_wysiwyg = "true";
defparam \regs[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[8]~483 (
// Equation(s):
// \rfif.rdat2[8]~483_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[25][8]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\regs[17][8]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[25][8]~q ),
	.datad(\regs[17][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~483_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~483 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[8]~483 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N21
dffeas \regs[21][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][8] .is_wysiwyg = "true";
defparam \regs[21][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N5
dffeas \regs[29][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][8] .is_wysiwyg = "true";
defparam \regs[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[8]~484 (
// Equation(s):
// \rfif.rdat2[8]~484_combout  = (Instr_IF_18 & ((\rfif.rdat2[8]~483_combout  & ((\regs[29][8]~q ))) # (!\rfif.rdat2[8]~483_combout  & (\regs[21][8]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[8]~483_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[8]~483_combout ),
	.datac(\regs[21][8]~q ),
	.datad(\regs[29][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~484_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~484 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[8]~484 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \regs[31][8]~feeder (
// Equation(s):
// \regs[31][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a6),
	.cin(gnd),
	.combout(\regs[31][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N9
dffeas \regs[31][8] (
	.clk(!CLK),
	.d(\regs[31][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][8] .is_wysiwyg = "true";
defparam \regs[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N27
dffeas \regs[19][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][8] .is_wysiwyg = "true";
defparam \regs[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \regs[27][8]~feeder (
// Equation(s):
// \regs[27][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a6),
	.cin(gnd),
	.combout(\regs[27][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \regs[27][8] (
	.clk(!CLK),
	.d(\regs[27][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][8] .is_wysiwyg = "true";
defparam \regs[27][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[8]~490 (
// Equation(s):
// \rfif.rdat2[8]~490_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[27][8]~q ))) # (!Instr_IF_19 & (\regs[19][8]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[19][8]~q ),
	.datad(\regs[27][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~490_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~490 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[8]~490 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[8]~491 (
// Equation(s):
// \rfif.rdat2[8]~491_combout  = (\rfif.rdat2[8]~490_combout  & (((\regs[31][8]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[8]~490_combout  & (\regs[23][8]~q  & ((Instr_IF_18))))

	.dataa(\regs[23][8]~q ),
	.datab(\regs[31][8]~q ),
	.datac(\rfif.rdat2[8]~490_combout ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~491_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~491 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[8]~491 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N3
dffeas \regs[30][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][8] .is_wysiwyg = "true";
defparam \regs[30][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N21
dffeas \regs[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][8] .is_wysiwyg = "true";
defparam \regs[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[8]~486 (
// Equation(s):
// \rfif.rdat2[8]~486_combout  = (\rfif.rdat2[8]~485_combout  & (((\regs[30][8]~q )) # (!Instr_IF_19))) # (!\rfif.rdat2[8]~485_combout  & (Instr_IF_19 & ((\regs[26][8]~q ))))

	.dataa(\rfif.rdat2[8]~485_combout ),
	.datab(Instr_IF_19),
	.datac(\regs[30][8]~q ),
	.datad(\regs[26][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~486_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~486 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[8]~486 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[8]~489 (
// Equation(s):
// \rfif.rdat2[8]~489_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[8]~486_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[8]~488_combout ))))

	.dataa(\rfif.rdat2[8]~488_combout ),
	.datab(Instr_IF_16),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[8]~486_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~489_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~489 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[8]~489 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \rfif.rdat2[8]~492 (
// Equation(s):
// \rfif.rdat2[8]~492_combout  = (\rfif.rdat2[8]~489_combout  & (((\rfif.rdat2[8]~491_combout ) # (!Instr_IF_16)))) # (!\rfif.rdat2[8]~489_combout  & (\rfif.rdat2[8]~484_combout  & ((Instr_IF_16))))

	.dataa(\rfif.rdat2[8]~484_combout ),
	.datab(\rfif.rdat2[8]~491_combout ),
	.datac(\rfif.rdat2[8]~489_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~492_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~492 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[8]~492 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \regs[7][8]~feeder (
// Equation(s):
// \regs[7][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[7][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[7][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N21
dffeas \regs[7][8] (
	.clk(!CLK),
	.d(\regs[7][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][8] .is_wysiwyg = "true";
defparam \regs[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N23
dffeas \regs[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][8] .is_wysiwyg = "true";
defparam \regs[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \regs[5][8]~feeder (
// Equation(s):
// \regs[5][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a6),
	.cin(gnd),
	.combout(\regs[5][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N13
dffeas \regs[5][8] (
	.clk(!CLK),
	.d(\regs[5][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][8] .is_wysiwyg = "true";
defparam \regs[5][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[8]~493 (
// Equation(s):
// \rfif.rdat2[8]~493_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[5][8]~q ))) # (!Instr_IF_16 & (\regs[4][8]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[4][8]~q ),
	.datad(\regs[5][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~493_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~493 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[8]~493 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \regs[6][8]~feeder (
// Equation(s):
// \regs[6][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a6),
	.cin(gnd),
	.combout(\regs[6][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[6][8]~feeder .lut_mask = 16'hFF00;
defparam \regs[6][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N19
dffeas \regs[6][8] (
	.clk(!CLK),
	.d(\regs[6][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][8] .is_wysiwyg = "true";
defparam \regs[6][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[8]~494 (
// Equation(s):
// \rfif.rdat2[8]~494_combout  = (Instr_IF_17 & ((\rfif.rdat2[8]~493_combout  & (\regs[7][8]~q )) # (!\rfif.rdat2[8]~493_combout  & ((\regs[6][8]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[8]~493_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[7][8]~q ),
	.datac(\rfif.rdat2[8]~493_combout ),
	.datad(\regs[6][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~494_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~494 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[8]~494 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \regs[15][8]~feeder (
// Equation(s):
// \regs[15][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N15
dffeas \regs[15][8] (
	.clk(!CLK),
	.d(\regs[15][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][8] .is_wysiwyg = "true";
defparam \regs[15][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N15
dffeas \regs[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][8] .is_wysiwyg = "true";
defparam \regs[12][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N1
dffeas \regs[13][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][8] .is_wysiwyg = "true";
defparam \regs[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \rfif.rdat2[8]~500 (
// Equation(s):
// \rfif.rdat2[8]~500_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][8]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][8]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][8]~q ),
	.datad(\regs[13][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~500_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~500 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[8]~500 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \regs[14][8]~feeder (
// Equation(s):
// \regs[14][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[14][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N21
dffeas \regs[14][8] (
	.clk(!CLK),
	.d(\regs[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][8] .is_wysiwyg = "true";
defparam \regs[14][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \rfif.rdat2[8]~501 (
// Equation(s):
// \rfif.rdat2[8]~501_combout  = (Instr_IF_17 & ((\rfif.rdat2[8]~500_combout  & (\regs[15][8]~q )) # (!\rfif.rdat2[8]~500_combout  & ((\regs[14][8]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[8]~500_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[15][8]~q ),
	.datac(\rfif.rdat2[8]~500_combout ),
	.datad(\regs[14][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~501_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~501 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[8]~501 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N17
dffeas \regs[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][8] .is_wysiwyg = "true";
defparam \regs[1][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N19
dffeas \regs[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][8] .is_wysiwyg = "true";
defparam \regs[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N27
dffeas \regs[0][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][8] .is_wysiwyg = "true";
defparam \regs[0][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \regs[2][8]~feeder (
// Equation(s):
// \regs[2][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N25
dffeas \regs[2][8] (
	.clk(!CLK),
	.d(\regs[2][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][8] .is_wysiwyg = "true";
defparam \regs[2][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[8]~497 (
// Equation(s):
// \rfif.rdat2[8]~497_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][8]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][8]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][8]~q ),
	.datad(\regs[2][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~497_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~497 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[8]~497 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[8]~498 (
// Equation(s):
// \rfif.rdat2[8]~498_combout  = (Instr_IF_16 & ((\rfif.rdat2[8]~497_combout  & ((\regs[3][8]~q ))) # (!\rfif.rdat2[8]~497_combout  & (\regs[1][8]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[8]~497_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][8]~q ),
	.datac(\regs[3][8]~q ),
	.datad(\rfif.rdat2[8]~497_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~498_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~498 .lut_mask = 16'hF588;
defparam \rfif.rdat2[8]~498 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N9
dffeas \regs[9][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][8] .is_wysiwyg = "true";
defparam \regs[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N11
dffeas \regs[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][8] .is_wysiwyg = "true";
defparam \regs[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N5
dffeas \regs[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][8] .is_wysiwyg = "true";
defparam \regs[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \regs[8][8]~feeder (
// Equation(s):
// \regs[8][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N3
dffeas \regs[8][8] (
	.clk(!CLK),
	.d(\regs[8][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][8] .is_wysiwyg = "true";
defparam \regs[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \rfif.rdat2[8]~495 (
// Equation(s):
// \rfif.rdat2[8]~495_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[10][8]~q )) # (!Instr_IF_17 & ((\regs[8][8]~q )))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[10][8]~q ),
	.datad(\regs[8][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~495_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~495 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[8]~495 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \rfif.rdat2[8]~496 (
// Equation(s):
// \rfif.rdat2[8]~496_combout  = (Instr_IF_16 & ((\rfif.rdat2[8]~495_combout  & ((\regs[11][8]~q ))) # (!\rfif.rdat2[8]~495_combout  & (\regs[9][8]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[8]~495_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[9][8]~q ),
	.datac(\regs[11][8]~q ),
	.datad(\rfif.rdat2[8]~495_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~496_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~496 .lut_mask = 16'hF588;
defparam \rfif.rdat2[8]~496 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \rfif.rdat2[8]~499 (
// Equation(s):
// \rfif.rdat2[8]~499_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\rfif.rdat2[8]~496_combout ))) # (!Instr_IF_19 & (\rfif.rdat2[8]~498_combout ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[8]~498_combout ),
	.datad(\rfif.rdat2[8]~496_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~499_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~499 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[8]~499 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[8]~502 (
// Equation(s):
// \rfif.rdat2[8]~502_combout  = (Instr_IF_18 & ((\rfif.rdat2[8]~499_combout  & ((\rfif.rdat2[8]~501_combout ))) # (!\rfif.rdat2[8]~499_combout  & (\rfif.rdat2[8]~494_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[8]~499_combout ))))

	.dataa(\rfif.rdat2[8]~494_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[8]~501_combout ),
	.datad(\rfif.rdat2[8]~499_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[8]~502_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[8]~502 .lut_mask = 16'hF388;
defparam \rfif.rdat2[8]~502 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N31
dffeas \regs[18][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][8] .is_wysiwyg = "true";
defparam \regs[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[8]~460 (
// Equation(s):
// \rfif.rdat1[8]~460_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][8]~q )) # (!Instr_IF_24 & ((\regs[18][8]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][8]~q ),
	.datad(\regs[18][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~460_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~460 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[8]~460 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N17
dffeas \regs[22][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][8] .is_wysiwyg = "true";
defparam \regs[22][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[8]~461 (
// Equation(s):
// \rfif.rdat1[8]~461_combout  = (\rfif.rdat1[8]~460_combout  & ((\regs[30][8]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[8]~460_combout  & (((\regs[22][8]~q  & Instr_IF_23))))

	.dataa(\regs[30][8]~q ),
	.datab(\rfif.rdat1[8]~460_combout ),
	.datac(\regs[22][8]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~461_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~461 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[8]~461 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \rfif.rdat1[8]~462 (
// Equation(s):
// \rfif.rdat1[8]~462_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][8]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[17][8]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[17][8]~q ),
	.datad(\regs[21][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~462_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~462 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[8]~462 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[8]~463 (
// Equation(s):
// \rfif.rdat1[8]~463_combout  = (Instr_IF_24 & ((\rfif.rdat1[8]~462_combout  & ((\regs[29][8]~q ))) # (!\rfif.rdat1[8]~462_combout  & (\regs[25][8]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[8]~462_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[25][8]~q ),
	.datac(\regs[29][8]~q ),
	.datad(\rfif.rdat1[8]~462_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~463_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~463 .lut_mask = 16'hF588;
defparam \rfif.rdat1[8]~463 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \regs[28][8]~feeder (
// Equation(s):
// \regs[28][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N23
dffeas \regs[28][8] (
	.clk(!CLK),
	.d(\regs[28][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][8] .is_wysiwyg = "true";
defparam \regs[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \regs[20][8]~feeder (
// Equation(s):
// \regs[20][8]~feeder_combout  = \input_a~111_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a6),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][8]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N29
dffeas \regs[20][8] (
	.clk(!CLK),
	.d(\regs[20][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][8] .is_wysiwyg = "true";
defparam \regs[20][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[8]~465 (
// Equation(s):
// \rfif.rdat1[8]~465_combout  = (\rfif.rdat1[8]~464_combout  & (((\regs[28][8]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[8]~464_combout  & (Instr_IF_23 & ((\regs[20][8]~q ))))

	.dataa(\rfif.rdat1[8]~464_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[28][8]~q ),
	.datad(\regs[20][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~465_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~465 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[8]~465 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \rfif.rdat1[8]~466 (
// Equation(s):
// \rfif.rdat1[8]~466_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\rfif.rdat1[8]~463_combout )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\rfif.rdat1[8]~465_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[8]~463_combout ),
	.datad(\rfif.rdat1[8]~465_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~466_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~466 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[8]~466 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N7
dffeas \regs[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][8] .is_wysiwyg = "true";
defparam \regs[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N6
cycloneive_lcell_comb \rfif.rdat1[8]~467 (
// Equation(s):
// \rfif.rdat1[8]~467_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[23][8]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & ((\regs[19][8]~q ))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[23][8]~q ),
	.datad(\regs[19][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~467_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~467 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[8]~467 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[8]~468 (
// Equation(s):
// \rfif.rdat1[8]~468_combout  = (\rfif.rdat1[8]~467_combout  & (((\regs[31][8]~q ) # (!Instr_IF_24)))) # (!\rfif.rdat1[8]~467_combout  & (\regs[27][8]~q  & ((Instr_IF_24))))

	.dataa(\rfif.rdat1[8]~467_combout ),
	.datab(\regs[27][8]~q ),
	.datac(\regs[31][8]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~468_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~468 .lut_mask = 16'hE4AA;
defparam \rfif.rdat1[8]~468 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \rfif.rdat1[8]~470 (
// Equation(s):
// \rfif.rdat1[8]~470_combout  = (Instr_IF_21 & (((\regs[9][8]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[8][8]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[8][8]~q ),
	.datac(\regs[9][8]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~470_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~470 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[8]~470 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \rfif.rdat1[8]~471 (
// Equation(s):
// \rfif.rdat1[8]~471_combout  = (Instr_IF_22 & ((\rfif.rdat1[8]~470_combout  & (\regs[11][8]~q )) # (!\rfif.rdat1[8]~470_combout  & ((\regs[10][8]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[8]~470_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[11][8]~q ),
	.datac(\regs[10][8]~q ),
	.datad(\rfif.rdat1[8]~470_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~471_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~471 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[8]~471 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \rfif.rdat1[8]~477 (
// Equation(s):
// \rfif.rdat1[8]~477_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][8]~q )) # (!Instr_IF_22 & ((\regs[12][8]~q )))))

	.dataa(Instr_IF_21),
	.datab(\regs[14][8]~q ),
	.datac(\regs[12][8]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~477_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~477 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[8]~477 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \rfif.rdat1[8]~478 (
// Equation(s):
// \rfif.rdat1[8]~478_combout  = (Instr_IF_21 & ((\rfif.rdat1[8]~477_combout  & (\regs[15][8]~q )) # (!\rfif.rdat1[8]~477_combout  & ((\regs[13][8]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[8]~477_combout ))))

	.dataa(\regs[15][8]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][8]~q ),
	.datad(\rfif.rdat1[8]~477_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~478_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~478 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[8]~478 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \rfif.rdat1[8]~472 (
// Equation(s):
// \rfif.rdat1[8]~472_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[6][8]~q ))) # (!Instr_IF_22 & (\regs[4][8]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[4][8]~q ),
	.datad(\regs[6][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~472_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~472 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[8]~472 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[8]~473 (
// Equation(s):
// \rfif.rdat1[8]~473_combout  = (Instr_IF_21 & ((\rfif.rdat1[8]~472_combout  & ((\regs[7][8]~q ))) # (!\rfif.rdat1[8]~472_combout  & (\regs[5][8]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[8]~472_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[5][8]~q ),
	.datac(\rfif.rdat1[8]~472_combout ),
	.datad(\regs[7][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~473_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~473 .lut_mask = 16'hF858;
defparam \rfif.rdat1[8]~473 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[8]~474 (
// Equation(s):
// \rfif.rdat1[8]~474_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][8]~q )) # (!Instr_IF_21 & ((\regs[0][8]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][8]~q ),
	.datad(\regs[0][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~474_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~474 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[8]~474 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[8]~475 (
// Equation(s):
// \rfif.rdat1[8]~475_combout  = (Instr_IF_22 & ((\rfif.rdat1[8]~474_combout  & (\regs[3][8]~q )) # (!\rfif.rdat1[8]~474_combout  & ((\regs[2][8]~q ))))) # (!Instr_IF_22 & (\rfif.rdat1[8]~474_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[8]~474_combout ),
	.datac(\regs[3][8]~q ),
	.datad(\regs[2][8]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~475_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~475 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[8]~475 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[8]~476 (
// Equation(s):
// \rfif.rdat1[8]~476_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & (\rfif.rdat1[8]~473_combout )) # (!Instr_IF_23 & ((\rfif.rdat1[8]~475_combout )))))

	.dataa(\rfif.rdat1[8]~473_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[8]~475_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[8]~476_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[8]~476 .lut_mask = 16'hEE30;
defparam \rfif.rdat1[8]~476 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N7
dffeas \regs[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][7] .is_wysiwyg = "true";
defparam \regs[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N30
cycloneive_lcell_comb \regs[9][7]~feeder (
// Equation(s):
// \regs[9][7]~feeder_combout  = \input_a~114_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][7]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N31
dffeas \regs[9][7] (
	.clk(!CLK),
	.d(\regs[9][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][7] .is_wysiwyg = "true";
defparam \regs[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[7]~514 (
// Equation(s):
// \rfif.rdat2[7]~514_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][7]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][7]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][7]~q ),
	.datad(\regs[9][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~514_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~514 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[7]~514 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N9
dffeas \regs[11][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][7] .is_wysiwyg = "true";
defparam \regs[11][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N8
cycloneive_lcell_comb \rfif.rdat2[7]~515 (
// Equation(s):
// \rfif.rdat2[7]~515_combout  = (\rfif.rdat2[7]~514_combout  & (((\regs[11][7]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[7]~514_combout  & (\regs[10][7]~q  & ((Instr_IF_17))))

	.dataa(\regs[10][7]~q ),
	.datab(\rfif.rdat2[7]~514_combout ),
	.datac(\regs[11][7]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~515_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~515 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[7]~515 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N5
dffeas \regs[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][7] .is_wysiwyg = "true";
defparam \regs[12][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N17
dffeas \regs[14][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][7] .is_wysiwyg = "true";
defparam \regs[14][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \rfif.rdat2[7]~521 (
// Equation(s):
// \rfif.rdat2[7]~521_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[14][7]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[12][7]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][7]~q ),
	.datad(\regs[14][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~521_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~521 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[7]~521 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \regs[13][7]~feeder (
// Equation(s):
// \regs[13][7]~feeder_combout  = \input_a~114_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][7]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N11
dffeas \regs[13][7] (
	.clk(!CLK),
	.d(\regs[13][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][7] .is_wysiwyg = "true";
defparam \regs[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N23
dffeas \regs[15][7] (
	.clk(!CLK),
	.d(input_a7),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][7] .is_wysiwyg = "true";
defparam \regs[15][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \rfif.rdat2[7]~522 (
// Equation(s):
// \rfif.rdat2[7]~522_combout  = (Instr_IF_16 & ((\rfif.rdat2[7]~521_combout  & ((\regs[15][7]~q ))) # (!\rfif.rdat2[7]~521_combout  & (\regs[13][7]~q )))) # (!Instr_IF_16 & (\rfif.rdat2[7]~521_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[7]~521_combout ),
	.datac(\regs[13][7]~q ),
	.datad(\regs[15][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~522_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~522 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[7]~522 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N19
dffeas \regs[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][7] .is_wysiwyg = "true";
defparam \regs[4][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N17
dffeas \regs[6][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][7] .is_wysiwyg = "true";
defparam \regs[6][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \rfif.rdat2[7]~516 (
// Equation(s):
// \rfif.rdat2[7]~516_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][7]~q ))) # (!Instr_IF_17 & (\regs[4][7]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][7]~q ),
	.datad(\regs[6][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~516_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~516 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[7]~516 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N19
dffeas \regs[7][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][7] .is_wysiwyg = "true";
defparam \regs[7][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N1
dffeas \regs[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][7] .is_wysiwyg = "true";
defparam \regs[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \rfif.rdat2[7]~517 (
// Equation(s):
// \rfif.rdat2[7]~517_combout  = (Instr_IF_16 & ((\rfif.rdat2[7]~516_combout  & (\regs[7][7]~q )) # (!\rfif.rdat2[7]~516_combout  & ((\regs[5][7]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[7]~516_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[7]~516_combout ),
	.datac(\regs[7][7]~q ),
	.datad(\regs[5][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~517_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~517 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[7]~517 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \regs[3][7]~feeder (
// Equation(s):
// \regs[3][7]~feeder_combout  = \input_a~114_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a7),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[3][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[3][7]~feeder .lut_mask = 16'hF0F0;
defparam \regs[3][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N17
dffeas \regs[3][7] (
	.clk(!CLK),
	.d(\regs[3][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][7] .is_wysiwyg = "true";
defparam \regs[3][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N1
dffeas \regs[2][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][7] .is_wysiwyg = "true";
defparam \regs[2][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N11
dffeas \regs[0][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][7] .is_wysiwyg = "true";
defparam \regs[0][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N31
dffeas \regs[1][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][7] .is_wysiwyg = "true";
defparam \regs[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[7]~518 (
// Equation(s):
// \rfif.rdat2[7]~518_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][7]~q ))) # (!Instr_IF_16 & (\regs[0][7]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][7]~q ),
	.datad(\regs[1][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~518_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~518 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[7]~518 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \rfif.rdat2[7]~519 (
// Equation(s):
// \rfif.rdat2[7]~519_combout  = (Instr_IF_17 & ((\rfif.rdat2[7]~518_combout  & (\regs[3][7]~q )) # (!\rfif.rdat2[7]~518_combout  & ((\regs[2][7]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[7]~518_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[3][7]~q ),
	.datac(\regs[2][7]~q ),
	.datad(\rfif.rdat2[7]~518_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~519_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~519 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[7]~519 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \rfif.rdat2[7]~520 (
// Equation(s):
// \rfif.rdat2[7]~520_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\rfif.rdat2[7]~517_combout )))) # (!Instr_IF_18 & (!Instr_IF_19 & ((\rfif.rdat2[7]~519_combout ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[7]~517_combout ),
	.datad(\rfif.rdat2[7]~519_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~520_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~520 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[7]~520 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[7]~523 (
// Equation(s):
// \rfif.rdat2[7]~523_combout  = (Instr_IF_19 & ((\rfif.rdat2[7]~520_combout  & ((\rfif.rdat2[7]~522_combout ))) # (!\rfif.rdat2[7]~520_combout  & (\rfif.rdat2[7]~515_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[7]~520_combout ))))

	.dataa(\rfif.rdat2[7]~515_combout ),
	.datab(\rfif.rdat2[7]~522_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[7]~520_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~523_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~523 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[7]~523 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N21
dffeas \regs[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][7] .is_wysiwyg = "true";
defparam \regs[22][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N27
dffeas \regs[18][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][7] .is_wysiwyg = "true";
defparam \regs[18][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N21
dffeas \regs[26][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][7] .is_wysiwyg = "true";
defparam \regs[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[7]~504 (
// Equation(s):
// \rfif.rdat2[7]~504_combout  = (Instr_IF_19 & (((\regs[26][7]~q ) # (Instr_IF_18)))) # (!Instr_IF_19 & (\regs[18][7]~q  & ((!Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[18][7]~q ),
	.datac(\regs[26][7]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~504_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~504 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[7]~504 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[7]~505 (
// Equation(s):
// \rfif.rdat2[7]~505_combout  = (Instr_IF_18 & ((\rfif.rdat2[7]~504_combout  & (\regs[30][7]~q )) # (!\rfif.rdat2[7]~504_combout  & ((\regs[22][7]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[7]~504_combout ))))

	.dataa(\regs[30][7]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][7]~q ),
	.datad(\rfif.rdat2[7]~504_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~505_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~505 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[7]~505 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \regs[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][7] .is_wysiwyg = "true";
defparam \regs[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \regs[23][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][7] .is_wysiwyg = "true";
defparam \regs[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[7]~511 (
// Equation(s):
// \rfif.rdat2[7]~511_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[23][7]~q ))) # (!Instr_IF_18 & (\regs[19][7]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[19][7]~q ),
	.datad(\regs[23][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~511_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~511 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[7]~511 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N11
dffeas \regs[31][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][7] .is_wysiwyg = "true";
defparam \regs[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N17
dffeas \regs[27][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][7] .is_wysiwyg = "true";
defparam \regs[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[7]~512 (
// Equation(s):
// \rfif.rdat2[7]~512_combout  = (Instr_IF_19 & ((\rfif.rdat2[7]~511_combout  & (\regs[31][7]~q )) # (!\rfif.rdat2[7]~511_combout  & ((\regs[27][7]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[7]~511_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[7]~511_combout ),
	.datac(\regs[31][7]~q ),
	.datad(\regs[27][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~512_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~512 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[7]~512 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N9
dffeas \regs[25][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][7] .is_wysiwyg = "true";
defparam \regs[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N31
dffeas \regs[29][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][7] .is_wysiwyg = "true";
defparam \regs[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N7
dffeas \regs[17][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][7] .is_wysiwyg = "true";
defparam \regs[17][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N25
dffeas \regs[21][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][7] .is_wysiwyg = "true";
defparam \regs[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N6
cycloneive_lcell_comb \rfif.rdat2[7]~506 (
// Equation(s):
// \rfif.rdat2[7]~506_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][7]~q ))) # (!Instr_IF_18 & (\regs[17][7]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][7]~q ),
	.datad(\regs[21][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~506_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~506 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[7]~506 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \rfif.rdat2[7]~507 (
// Equation(s):
// \rfif.rdat2[7]~507_combout  = (Instr_IF_19 & ((\rfif.rdat2[7]~506_combout  & ((\regs[29][7]~q ))) # (!\rfif.rdat2[7]~506_combout  & (\regs[25][7]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[7]~506_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][7]~q ),
	.datac(\regs[29][7]~q ),
	.datad(\rfif.rdat2[7]~506_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~507_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~507 .lut_mask = 16'hF588;
defparam \rfif.rdat2[7]~507 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \rfif.rdat2[7]~510 (
// Equation(s):
// \rfif.rdat2[7]~510_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\rfif.rdat2[7]~507_combout ))) # (!Instr_IF_16 & (\rfif.rdat2[7]~509_combout ))))

	.dataa(\rfif.rdat2[7]~509_combout ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[7]~507_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~510_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~510 .lut_mask = 16'hF2C2;
defparam \rfif.rdat2[7]~510 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[7]~513 (
// Equation(s):
// \rfif.rdat2[7]~513_combout  = (Instr_IF_17 & ((\rfif.rdat2[7]~510_combout  & ((\rfif.rdat2[7]~512_combout ))) # (!\rfif.rdat2[7]~510_combout  & (\rfif.rdat2[7]~505_combout )))) # (!Instr_IF_17 & (((\rfif.rdat2[7]~510_combout ))))

	.dataa(\rfif.rdat2[7]~505_combout ),
	.datab(\rfif.rdat2[7]~512_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[7]~510_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[7]~513_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[7]~513 .lut_mask = 16'hCFA0;
defparam \rfif.rdat2[7]~513 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \rfif.rdat1[7]~480 (
// Equation(s):
// \rfif.rdat1[7]~480_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][7]~q ))) # (!Instr_IF_24 & (\regs[17][7]~q ))))

	.dataa(\regs[17][7]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[25][7]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~480_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~480 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[7]~480 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[7]~481 (
// Equation(s):
// \rfif.rdat1[7]~481_combout  = (Instr_IF_23 & ((\rfif.rdat1[7]~480_combout  & (\regs[29][7]~q )) # (!\rfif.rdat1[7]~480_combout  & ((\regs[21][7]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[7]~480_combout ))))

	.dataa(\regs[29][7]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[21][7]~q ),
	.datad(\rfif.rdat1[7]~480_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~481_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~481 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[7]~481 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[7]~487 (
// Equation(s):
// \rfif.rdat1[7]~487_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][7]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][7]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][7]~q ),
	.datad(\regs[19][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~487_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~487 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[7]~487 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[7]~488 (
// Equation(s):
// \rfif.rdat1[7]~488_combout  = (Instr_IF_23 & ((\rfif.rdat1[7]~487_combout  & (\regs[31][7]~q )) # (!\rfif.rdat1[7]~487_combout  & ((\regs[23][7]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[7]~487_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[31][7]~q ),
	.datac(\regs[23][7]~q ),
	.datad(\rfif.rdat1[7]~487_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~488_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~488 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[7]~488 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N5
dffeas \regs[20][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][7] .is_wysiwyg = "true";
defparam \regs[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[7]~484 (
// Equation(s):
// \rfif.rdat1[7]~484_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[20][7]~q ))) # (!Instr_IF_23 & (\regs[16][7]~q ))))

	.dataa(\regs[16][7]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[20][7]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~484_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~484 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[7]~484 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N5
dffeas \regs[24][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][7] .is_wysiwyg = "true";
defparam \regs[24][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[7]~485 (
// Equation(s):
// \rfif.rdat1[7]~485_combout  = (\rfif.rdat1[7]~484_combout  & ((\regs[28][7]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[7]~484_combout  & (((\regs[24][7]~q  & Instr_IF_24))))

	.dataa(\regs[28][7]~q ),
	.datab(\rfif.rdat1[7]~484_combout ),
	.datac(\regs[24][7]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~485_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~485 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[7]~485 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \rfif.rdat1[7]~482 (
// Equation(s):
// \rfif.rdat1[7]~482_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][7]~q ))) # (!Instr_IF_23 & (\regs[18][7]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[18][7]~q ),
	.datad(\regs[22][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~482_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~482 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[7]~482 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N15
dffeas \regs[30][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][7] .is_wysiwyg = "true";
defparam \regs[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \rfif.rdat1[7]~483 (
// Equation(s):
// \rfif.rdat1[7]~483_combout  = (Instr_IF_24 & ((\rfif.rdat1[7]~482_combout  & (\regs[30][7]~q )) # (!\rfif.rdat1[7]~482_combout  & ((\regs[26][7]~q ))))) # (!Instr_IF_24 & (\rfif.rdat1[7]~482_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[7]~482_combout ),
	.datac(\regs[30][7]~q ),
	.datad(\regs[26][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~483_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~483 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[7]~483 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \rfif.rdat1[7]~486 (
// Equation(s):
// \rfif.rdat1[7]~486_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\rfif.rdat1[7]~483_combout ))) # (!Instr_IF_22 & (\rfif.rdat1[7]~485_combout ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[7]~485_combout ),
	.datad(\rfif.rdat1[7]~483_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~486_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~486 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[7]~486 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N17
dffeas \regs[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][7] .is_wysiwyg = "true";
defparam \regs[10][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[7]~492 (
// Equation(s):
// \rfif.rdat1[7]~492_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][7]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][7]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][7]~q ),
	.datad(\regs[8][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~492_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~492 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[7]~492 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N18
cycloneive_lcell_comb \rfif.rdat1[7]~493 (
// Equation(s):
// \rfif.rdat1[7]~493_combout  = (Instr_IF_21 & ((\rfif.rdat1[7]~492_combout  & (\regs[11][7]~q )) # (!\rfif.rdat1[7]~492_combout  & ((\regs[9][7]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[7]~492_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[11][7]~q ),
	.datac(\regs[9][7]~q ),
	.datad(\rfif.rdat1[7]~492_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~493_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~493 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[7]~493 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[7]~494 (
// Equation(s):
// \rfif.rdat1[7]~494_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[2][7]~q ))) # (!Instr_IF_22 & (\regs[0][7]~q ))))

	.dataa(Instr_IF_21),
	.datab(\regs[0][7]~q ),
	.datac(Instr_IF_22),
	.datad(\regs[2][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~494_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~494 .lut_mask = 16'hF4A4;
defparam \rfif.rdat1[7]~494 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \rfif.rdat1[7]~495 (
// Equation(s):
// \rfif.rdat1[7]~495_combout  = (Instr_IF_21 & ((\rfif.rdat1[7]~494_combout  & ((\regs[3][7]~q ))) # (!\rfif.rdat1[7]~494_combout  & (\regs[1][7]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[7]~494_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[7]~494_combout ),
	.datac(\regs[1][7]~q ),
	.datad(\regs[3][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~495_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~495 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[7]~495 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \rfif.rdat1[7]~496 (
// Equation(s):
// \rfif.rdat1[7]~496_combout  = (Instr_IF_24 & ((\rfif.rdat1[7]~493_combout ) # ((Instr_IF_23)))) # (!Instr_IF_24 & (((\rfif.rdat1[7]~495_combout  & !Instr_IF_23))))

	.dataa(\rfif.rdat1[7]~493_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[7]~495_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~496_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~496 .lut_mask = 16'hCCB8;
defparam \rfif.rdat1[7]~496 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[7]~490 (
// Equation(s):
// \rfif.rdat1[7]~490_combout  = (Instr_IF_21 & (((\regs[5][7]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[4][7]~q  & ((!Instr_IF_22))))

	.dataa(\regs[4][7]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][7]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~490_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~490 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[7]~490 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \rfif.rdat1[7]~491 (
// Equation(s):
// \rfif.rdat1[7]~491_combout  = (\rfif.rdat1[7]~490_combout  & ((\regs[7][7]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[7]~490_combout  & (((\regs[6][7]~q  & Instr_IF_22))))

	.dataa(\rfif.rdat1[7]~490_combout ),
	.datab(\regs[7][7]~q ),
	.datac(\regs[6][7]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~491_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~491 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[7]~491 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \rfif.rdat1[7]~497 (
// Equation(s):
// \rfif.rdat1[7]~497_combout  = (Instr_IF_21 & ((\regs[13][7]~q ) # ((Instr_IF_22)))) # (!Instr_IF_21 & (((!Instr_IF_22 & \regs[12][7]~q ))))

	.dataa(\regs[13][7]~q ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\regs[12][7]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~497_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~497 .lut_mask = 16'hCBC8;
defparam \rfif.rdat1[7]~497 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \rfif.rdat1[7]~498 (
// Equation(s):
// \rfif.rdat1[7]~498_combout  = (Instr_IF_22 & ((\rfif.rdat1[7]~497_combout  & (\regs[15][7]~q )) # (!\rfif.rdat1[7]~497_combout  & ((\regs[14][7]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[7]~497_combout ))))

	.dataa(\regs[15][7]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[14][7]~q ),
	.datad(\rfif.rdat1[7]~497_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[7]~498_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[7]~498 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[7]~498 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N5
dffeas \regs[26][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][6] .is_wysiwyg = "true";
defparam \regs[26][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N31
dffeas \regs[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][6] .is_wysiwyg = "true";
defparam \regs[30][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N9
dffeas \regs[22][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][6] .is_wysiwyg = "true";
defparam \regs[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N27
dffeas \regs[18][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][6] .is_wysiwyg = "true";
defparam \regs[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[6]~527 (
// Equation(s):
// \rfif.rdat2[6]~527_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[22][6]~q )) # (!Instr_IF_18 & ((\regs[18][6]~q )))))

	.dataa(Instr_IF_19),
	.datab(\regs[22][6]~q ),
	.datac(\regs[18][6]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~527_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~527 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[6]~527 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \rfif.rdat2[6]~528 (
// Equation(s):
// \rfif.rdat2[6]~528_combout  = (Instr_IF_19 & ((\rfif.rdat2[6]~527_combout  & ((\regs[30][6]~q ))) # (!\rfif.rdat2[6]~527_combout  & (\regs[26][6]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[6]~527_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][6]~q ),
	.datac(\regs[30][6]~q ),
	.datad(\rfif.rdat2[6]~527_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~528_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~528 .lut_mask = 16'hF588;
defparam \rfif.rdat2[6]~528 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[6]~531 (
// Equation(s):
// \rfif.rdat2[6]~531_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[6]~528_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[6]~530_combout ))))

	.dataa(\rfif.rdat2[6]~530_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[6]~528_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~531_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~531 .lut_mask = 16'hFC22;
defparam \rfif.rdat2[6]~531 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N29
dffeas \regs[21][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][6] .is_wysiwyg = "true";
defparam \regs[21][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N19
dffeas \regs[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][6] .is_wysiwyg = "true";
defparam \regs[17][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N27
dffeas \regs[25][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][6] .is_wysiwyg = "true";
defparam \regs[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[6]~525 (
// Equation(s):
// \rfif.rdat2[6]~525_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][6]~q ))) # (!Instr_IF_19 & (\regs[17][6]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[17][6]~q ),
	.datac(\regs[25][6]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~525_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~525 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[6]~525 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \rfif.rdat2[6]~526 (
// Equation(s):
// \rfif.rdat2[6]~526_combout  = (Instr_IF_18 & ((\rfif.rdat2[6]~525_combout  & (\regs[29][6]~q )) # (!\rfif.rdat2[6]~525_combout  & ((\regs[21][6]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[6]~525_combout ))))

	.dataa(\regs[29][6]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[21][6]~q ),
	.datad(\rfif.rdat2[6]~525_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~526_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~526 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[6]~526 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N21
dffeas \regs[23][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][6] .is_wysiwyg = "true";
defparam \regs[23][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \regs[31][6]~feeder (
// Equation(s):
// \regs[31][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a8),
	.cin(gnd),
	.combout(\regs[31][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][6]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N5
dffeas \regs[31][6] (
	.clk(!CLK),
	.d(\regs[31][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][6] .is_wysiwyg = "true";
defparam \regs[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \rfif.rdat2[6]~533 (
// Equation(s):
// \rfif.rdat2[6]~533_combout  = (\rfif.rdat2[6]~532_combout  & (((\regs[31][6]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[6]~532_combout  & (\regs[23][6]~q  & ((Instr_IF_18))))

	.dataa(\rfif.rdat2[6]~532_combout ),
	.datab(\regs[23][6]~q ),
	.datac(\regs[31][6]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~533_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~533 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[6]~533 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[6]~534 (
// Equation(s):
// \rfif.rdat2[6]~534_combout  = (\rfif.rdat2[6]~531_combout  & (((\rfif.rdat2[6]~533_combout )) # (!Instr_IF_16))) # (!\rfif.rdat2[6]~531_combout  & (Instr_IF_16 & (\rfif.rdat2[6]~526_combout )))

	.dataa(\rfif.rdat2[6]~531_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[6]~526_combout ),
	.datad(\rfif.rdat2[6]~533_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~534_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~534 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[6]~534 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N17
dffeas \regs[6][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][6] .is_wysiwyg = "true";
defparam \regs[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N15
dffeas \regs[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][6] .is_wysiwyg = "true";
defparam \regs[5][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N11
dffeas \regs[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][6] .is_wysiwyg = "true";
defparam \regs[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[6]~535 (
// Equation(s):
// \rfif.rdat2[6]~535_combout  = (Instr_IF_16 & ((\regs[5][6]~q ) # ((Instr_IF_17)))) # (!Instr_IF_16 & (((\regs[4][6]~q  & !Instr_IF_17))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][6]~q ),
	.datac(\regs[4][6]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~535_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~535 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[6]~535 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \rfif.rdat2[6]~536 (
// Equation(s):
// \rfif.rdat2[6]~536_combout  = (Instr_IF_17 & ((\rfif.rdat2[6]~535_combout  & (\regs[7][6]~q )) # (!\rfif.rdat2[6]~535_combout  & ((\regs[6][6]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[6]~535_combout ))))

	.dataa(\regs[7][6]~q ),
	.datab(\regs[6][6]~q ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[6]~535_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~536_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~536 .lut_mask = 16'hAFC0;
defparam \rfif.rdat2[6]~536 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \regs[15][6]~feeder (
// Equation(s):
// \regs[15][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[15][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[15][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \regs[15][6] (
	.clk(!CLK),
	.d(\regs[15][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][6] .is_wysiwyg = "true";
defparam \regs[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N27
dffeas \regs[14][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][6] .is_wysiwyg = "true";
defparam \regs[14][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \rfif.rdat2[6]~543 (
// Equation(s):
// \rfif.rdat2[6]~543_combout  = (\rfif.rdat2[6]~542_combout  & ((\regs[15][6]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[6]~542_combout  & (((\regs[14][6]~q  & Instr_IF_17))))

	.dataa(\rfif.rdat2[6]~542_combout ),
	.datab(\regs[15][6]~q ),
	.datac(\regs[14][6]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~543_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~543 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[6]~543 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N17
dffeas \regs[1][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][6] .is_wysiwyg = "true";
defparam \regs[1][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N27
dffeas \regs[3][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][6] .is_wysiwyg = "true";
defparam \regs[3][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N17
dffeas \regs[0][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][6] .is_wysiwyg = "true";
defparam \regs[0][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \rfif.rdat2[6]~539 (
// Equation(s):
// \rfif.rdat2[6]~539_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][6]~q )) # (!Instr_IF_17 & ((\regs[0][6]~q )))))

	.dataa(\regs[2][6]~q ),
	.datab(Instr_IF_16),
	.datac(\regs[0][6]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~539_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~539 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[6]~539 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[6]~540 (
// Equation(s):
// \rfif.rdat2[6]~540_combout  = (Instr_IF_16 & ((\rfif.rdat2[6]~539_combout  & ((\regs[3][6]~q ))) # (!\rfif.rdat2[6]~539_combout  & (\regs[1][6]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[6]~539_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[1][6]~q ),
	.datac(\regs[3][6]~q ),
	.datad(\rfif.rdat2[6]~539_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~540_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~540 .lut_mask = 16'hF588;
defparam \rfif.rdat2[6]~540 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N31
dffeas \regs[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][6] .is_wysiwyg = "true";
defparam \regs[10][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N2
cycloneive_lcell_comb \regs[8][6]~feeder (
// Equation(s):
// \regs[8][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N3
dffeas \regs[8][6] (
	.clk(!CLK),
	.d(\regs[8][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][6] .is_wysiwyg = "true";
defparam \regs[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[6]~537 (
// Equation(s):
// \rfif.rdat2[6]~537_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[10][6]~q )) # (!Instr_IF_17 & ((\regs[8][6]~q )))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[10][6]~q ),
	.datad(\regs[8][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~537_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~537 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[6]~537 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N15
dffeas \regs[11][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][6] .is_wysiwyg = "true";
defparam \regs[11][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \regs[9][6]~feeder (
// Equation(s):
// \regs[9][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N13
dffeas \regs[9][6] (
	.clk(!CLK),
	.d(\regs[9][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][6] .is_wysiwyg = "true";
defparam \regs[9][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \rfif.rdat2[6]~538 (
// Equation(s):
// \rfif.rdat2[6]~538_combout  = (Instr_IF_16 & ((\rfif.rdat2[6]~537_combout  & (\regs[11][6]~q )) # (!\rfif.rdat2[6]~537_combout  & ((\regs[9][6]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[6]~537_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[6]~537_combout ),
	.datac(\regs[11][6]~q ),
	.datad(\regs[9][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~538_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~538 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[6]~538 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[6]~541 (
// Equation(s):
// \rfif.rdat2[6]~541_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\rfif.rdat2[6]~538_combout ))) # (!Instr_IF_19 & (\rfif.rdat2[6]~540_combout ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[6]~540_combout ),
	.datad(\rfif.rdat2[6]~538_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~541_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~541 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[6]~541 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \rfif.rdat2[6]~544 (
// Equation(s):
// \rfif.rdat2[6]~544_combout  = (Instr_IF_18 & ((\rfif.rdat2[6]~541_combout  & ((\rfif.rdat2[6]~543_combout ))) # (!\rfif.rdat2[6]~541_combout  & (\rfif.rdat2[6]~536_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[6]~541_combout ))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[6]~536_combout ),
	.datac(\rfif.rdat2[6]~543_combout ),
	.datad(\rfif.rdat2[6]~541_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[6]~544_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[6]~544 .lut_mask = 16'hF588;
defparam \rfif.rdat2[6]~544 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[6]~500 (
// Equation(s):
// \rfif.rdat1[6]~500_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][6]~q )) # (!Instr_IF_24 & ((\regs[18][6]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][6]~q ),
	.datad(\regs[18][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~500_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~500 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[6]~500 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[6]~501 (
// Equation(s):
// \rfif.rdat1[6]~501_combout  = (Instr_IF_23 & ((\rfif.rdat1[6]~500_combout  & ((\regs[30][6]~q ))) # (!\rfif.rdat1[6]~500_combout  & (\regs[22][6]~q )))) # (!Instr_IF_23 & (\rfif.rdat1[6]~500_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[6]~500_combout ),
	.datac(\regs[22][6]~q ),
	.datad(\regs[30][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~501_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~501 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[6]~501 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \regs[27][6]~feeder (
// Equation(s):
// \regs[27][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a8),
	.cin(gnd),
	.combout(\regs[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][6]~feeder .lut_mask = 16'hFF00;
defparam \regs[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N23
dffeas \regs[27][6] (
	.clk(!CLK),
	.d(\regs[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][6] .is_wysiwyg = "true";
defparam \regs[27][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N31
dffeas \regs[19][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][6] .is_wysiwyg = "true";
defparam \regs[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \rfif.rdat1[6]~507 (
// Equation(s):
// \rfif.rdat1[6]~507_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & (\regs[23][6]~q )) # (!Instr_IF_23 & ((\regs[19][6]~q )))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[23][6]~q ),
	.datad(\regs[19][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~507_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~507 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[6]~507 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[6]~508 (
// Equation(s):
// \rfif.rdat1[6]~508_combout  = (Instr_IF_24 & ((\rfif.rdat1[6]~507_combout  & (\regs[31][6]~q )) # (!\rfif.rdat1[6]~507_combout  & ((\regs[27][6]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[6]~507_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[31][6]~q ),
	.datac(\regs[27][6]~q ),
	.datad(\rfif.rdat1[6]~507_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~508_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~508 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[6]~508 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N4
cycloneive_lcell_comb \regs[20][6]~feeder (
// Equation(s):
// \regs[20][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[20][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[20][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N5
dffeas \regs[20][6] (
	.clk(!CLK),
	.d(\regs[20][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][6] .is_wysiwyg = "true";
defparam \regs[20][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \regs[28][6]~feeder (
// Equation(s):
// \regs[28][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[28][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[28][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N19
dffeas \regs[28][6] (
	.clk(!CLK),
	.d(\regs[28][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][6] .is_wysiwyg = "true";
defparam \regs[28][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \rfif.rdat1[6]~505 (
// Equation(s):
// \rfif.rdat1[6]~505_combout  = (\rfif.rdat1[6]~504_combout  & (((\regs[28][6]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[6]~504_combout  & (Instr_IF_23 & (\regs[20][6]~q )))

	.dataa(\rfif.rdat1[6]~504_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[20][6]~q ),
	.datad(\regs[28][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~505_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~505 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[6]~505 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[6]~502 (
// Equation(s):
// \rfif.rdat1[6]~502_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][6]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[17][6]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[17][6]~q ),
	.datad(\regs[21][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~502_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~502 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[6]~502 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N25
dffeas \regs[29][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][6] .is_wysiwyg = "true";
defparam \regs[29][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[6]~503 (
// Equation(s):
// \rfif.rdat1[6]~503_combout  = (\rfif.rdat1[6]~502_combout  & (((\regs[29][6]~q ) # (!Instr_IF_24)))) # (!\rfif.rdat1[6]~502_combout  & (\regs[25][6]~q  & ((Instr_IF_24))))

	.dataa(\regs[25][6]~q ),
	.datab(\rfif.rdat1[6]~502_combout ),
	.datac(\regs[29][6]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~503_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~503 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[6]~503 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[6]~506 (
// Equation(s):
// \rfif.rdat1[6]~506_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\rfif.rdat1[6]~503_combout ))) # (!Instr_IF_21 & (\rfif.rdat1[6]~505_combout ))))

	.dataa(\rfif.rdat1[6]~505_combout ),
	.datab(Instr_IF_22),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[6]~503_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~506_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~506 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[6]~506 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[6]~510 (
// Equation(s):
// \rfif.rdat1[6]~510_combout  = (Instr_IF_21 & ((\regs[9][6]~q ) # ((Instr_IF_22)))) # (!Instr_IF_21 & (((\regs[8][6]~q  & !Instr_IF_22))))

	.dataa(\regs[9][6]~q ),
	.datab(\regs[8][6]~q ),
	.datac(Instr_IF_21),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~510_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~510 .lut_mask = 16'hF0AC;
defparam \rfif.rdat1[6]~510 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[6]~511 (
// Equation(s):
// \rfif.rdat1[6]~511_combout  = (Instr_IF_22 & ((\rfif.rdat1[6]~510_combout  & ((\regs[11][6]~q ))) # (!\rfif.rdat1[6]~510_combout  & (\regs[10][6]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[6]~510_combout ))))

	.dataa(\regs[10][6]~q ),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[6]~510_combout ),
	.datad(\regs[11][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~511_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~511 .lut_mask = 16'hF838;
defparam \rfif.rdat1[6]~511 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \regs[2][6]~feeder (
// Equation(s):
// \regs[2][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N23
dffeas \regs[2][6] (
	.clk(!CLK),
	.d(\regs[2][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][6] .is_wysiwyg = "true";
defparam \regs[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \rfif.rdat1[6]~515 (
// Equation(s):
// \rfif.rdat1[6]~515_combout  = (\rfif.rdat1[6]~514_combout  & (((\regs[3][6]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[6]~514_combout  & (Instr_IF_22 & ((\regs[2][6]~q ))))

	.dataa(\rfif.rdat1[6]~514_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[3][6]~q ),
	.datad(\regs[2][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~515_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~515 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[6]~515 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \regs[7][6]~feeder (
// Equation(s):
// \regs[7][6]~feeder_combout  = \input_a~117_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a8),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[7][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][6]~feeder .lut_mask = 16'hF0F0;
defparam \regs[7][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N31
dffeas \regs[7][6] (
	.clk(!CLK),
	.d(\regs[7][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][6] .is_wysiwyg = "true";
defparam \regs[7][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[6]~513 (
// Equation(s):
// \rfif.rdat1[6]~513_combout  = (\rfif.rdat1[6]~512_combout  & (((\regs[7][6]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[6]~512_combout  & (Instr_IF_21 & (\regs[5][6]~q )))

	.dataa(\rfif.rdat1[6]~512_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[5][6]~q ),
	.datad(\regs[7][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~513_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~513 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[6]~513 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N16
cycloneive_lcell_comb \rfif.rdat1[6]~516 (
// Equation(s):
// \rfif.rdat1[6]~516_combout  = (Instr_IF_23 & (((\rfif.rdat1[6]~513_combout ) # (Instr_IF_24)))) # (!Instr_IF_23 & (\rfif.rdat1[6]~515_combout  & ((!Instr_IF_24))))

	.dataa(\rfif.rdat1[6]~515_combout ),
	.datab(\rfif.rdat1[6]~513_combout ),
	.datac(Instr_IF_23),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~516_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~516 .lut_mask = 16'hF0CA;
defparam \rfif.rdat1[6]~516 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N21
dffeas \regs[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][6] .is_wysiwyg = "true";
defparam \regs[13][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N27
dffeas \regs[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][6] .is_wysiwyg = "true";
defparam \regs[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[6]~517 (
// Equation(s):
// \rfif.rdat1[6]~517_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[14][6]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & (\regs[12][6]~q )))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[12][6]~q ),
	.datad(\regs[14][6]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~517_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~517 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[6]~517 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \rfif.rdat1[6]~518 (
// Equation(s):
// \rfif.rdat1[6]~518_combout  = (Instr_IF_21 & ((\rfif.rdat1[6]~517_combout  & (\regs[15][6]~q )) # (!\rfif.rdat1[6]~517_combout  & ((\regs[13][6]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[6]~517_combout ))))

	.dataa(\regs[15][6]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][6]~q ),
	.datad(\rfif.rdat1[6]~517_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[6]~518_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[6]~518 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[6]~518 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N15
dffeas \regs[28][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][5] .is_wysiwyg = "true";
defparam \regs[28][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N9
dffeas \regs[24][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][5] .is_wysiwyg = "true";
defparam \regs[24][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N15
dffeas \regs[16][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][5] .is_wysiwyg = "true";
defparam \regs[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[5]~550 (
// Equation(s):
// \rfif.rdat2[5]~550_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\regs[24][5]~q )) # (!Instr_IF_19 & ((\regs[16][5]~q )))))

	.dataa(Instr_IF_18),
	.datab(\regs[24][5]~q ),
	.datac(\regs[16][5]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~550_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~550 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[5]~550 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N14
cycloneive_lcell_comb \rfif.rdat2[5]~551 (
// Equation(s):
// \rfif.rdat2[5]~551_combout  = (Instr_IF_18 & ((\rfif.rdat2[5]~550_combout  & ((\regs[28][5]~q ))) # (!\rfif.rdat2[5]~550_combout  & (\regs[20][5]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[5]~550_combout ))))

	.dataa(\regs[20][5]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][5]~q ),
	.datad(\rfif.rdat2[5]~550_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~551_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~551 .lut_mask = 16'hF388;
defparam \rfif.rdat2[5]~551 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[5]~552 (
// Equation(s):
// \rfif.rdat2[5]~552_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[5]~549_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[5]~551_combout )))))

	.dataa(\rfif.rdat2[5]~549_combout ),
	.datab(Instr_IF_17),
	.datac(Instr_IF_16),
	.datad(\rfif.rdat2[5]~551_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~552_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~552 .lut_mask = 16'hE3E0;
defparam \rfif.rdat2[5]~552 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N21
dffeas \regs[27][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][5] .is_wysiwyg = "true";
defparam \regs[27][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N23
dffeas \regs[31][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][5] .is_wysiwyg = "true";
defparam \regs[31][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[5]~554 (
// Equation(s):
// \rfif.rdat2[5]~554_combout  = (\rfif.rdat2[5]~553_combout  & (((\regs[31][5]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[5]~553_combout  & (\regs[27][5]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[5]~553_combout ),
	.datab(\regs[27][5]~q ),
	.datac(\regs[31][5]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~554_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~554 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[5]~554 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N9
dffeas \regs[22][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][5] .is_wysiwyg = "true";
defparam \regs[22][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N23
dffeas \regs[30][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][5] .is_wysiwyg = "true";
defparam \regs[30][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \rfif.rdat2[5]~547 (
// Equation(s):
// \rfif.rdat2[5]~547_combout  = (\rfif.rdat2[5]~546_combout  & (((\regs[30][5]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[5]~546_combout  & (Instr_IF_18 & (\regs[22][5]~q )))

	.dataa(\rfif.rdat2[5]~546_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[22][5]~q ),
	.datad(\regs[30][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~547_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~547 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[5]~547 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[5]~555 (
// Equation(s):
// \rfif.rdat2[5]~555_combout  = (\rfif.rdat2[5]~552_combout  & ((\rfif.rdat2[5]~554_combout ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[5]~552_combout  & (((Instr_IF_17 & \rfif.rdat2[5]~547_combout ))))

	.dataa(\rfif.rdat2[5]~552_combout ),
	.datab(\rfif.rdat2[5]~554_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[5]~547_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~555_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~555 .lut_mask = 16'hDA8A;
defparam \rfif.rdat2[5]~555 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N5
dffeas \regs[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][5] .is_wysiwyg = "true";
defparam \regs[10][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N3
dffeas \regs[11][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][5] .is_wysiwyg = "true";
defparam \regs[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N11
dffeas \regs[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][5] .is_wysiwyg = "true";
defparam \regs[8][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N25
dffeas \regs[9][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][5] .is_wysiwyg = "true";
defparam \regs[9][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[5]~556 (
// Equation(s):
// \rfif.rdat2[5]~556_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[9][5]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[8][5]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[8][5]~q ),
	.datad(\regs[9][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~556_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~556 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[5]~556 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N2
cycloneive_lcell_comb \rfif.rdat2[5]~557 (
// Equation(s):
// \rfif.rdat2[5]~557_combout  = (Instr_IF_17 & ((\rfif.rdat2[5]~556_combout  & ((\regs[11][5]~q ))) # (!\rfif.rdat2[5]~556_combout  & (\regs[10][5]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[5]~556_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[10][5]~q ),
	.datac(\regs[11][5]~q ),
	.datad(\rfif.rdat2[5]~556_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~557_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~557 .lut_mask = 16'hF588;
defparam \rfif.rdat2[5]~557 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N20
cycloneive_lcell_comb \regs[12][5]~feeder (
// Equation(s):
// \regs[12][5]~feeder_combout  = \input_a~120_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a9),
	.cin(gnd),
	.combout(\regs[12][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[12][5]~feeder .lut_mask = 16'hFF00;
defparam \regs[12][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N21
dffeas \regs[12][5] (
	.clk(!CLK),
	.d(\regs[12][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][5] .is_wysiwyg = "true";
defparam \regs[12][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N29
dffeas \regs[14][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][5] .is_wysiwyg = "true";
defparam \regs[14][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[5]~563 (
// Equation(s):
// \rfif.rdat2[5]~563_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[14][5]~q ))) # (!Instr_IF_17 & (\regs[12][5]~q ))))

	.dataa(Instr_IF_16),
	.datab(\regs[12][5]~q ),
	.datac(Instr_IF_17),
	.datad(\regs[14][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~563_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~563 .lut_mask = 16'hF4A4;
defparam \rfif.rdat2[5]~563 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \regs[15][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][5] .is_wysiwyg = "true";
defparam \regs[15][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N2
cycloneive_lcell_comb \regs[13][5]~feeder (
// Equation(s):
// \regs[13][5]~feeder_combout  = \input_a~120_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a9),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[13][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[13][5]~feeder .lut_mask = 16'hF0F0;
defparam \regs[13][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N3
dffeas \regs[13][5] (
	.clk(!CLK),
	.d(\regs[13][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][5] .is_wysiwyg = "true";
defparam \regs[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[5]~564 (
// Equation(s):
// \rfif.rdat2[5]~564_combout  = (Instr_IF_16 & ((\rfif.rdat2[5]~563_combout  & (\regs[15][5]~q )) # (!\rfif.rdat2[5]~563_combout  & ((\regs[13][5]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[5]~563_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[5]~563_combout ),
	.datac(\regs[15][5]~q ),
	.datad(\regs[13][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~564_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~564 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[5]~564 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N21
dffeas \regs[2][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][5] .is_wysiwyg = "true";
defparam \regs[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N19
dffeas \regs[3][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][5] .is_wysiwyg = "true";
defparam \regs[3][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N3
dffeas \regs[0][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][5] .is_wysiwyg = "true";
defparam \regs[0][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N29
dffeas \regs[1][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][5] .is_wysiwyg = "true";
defparam \regs[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \rfif.rdat2[5]~560 (
// Equation(s):
// \rfif.rdat2[5]~560_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[1][5]~q ))) # (!Instr_IF_16 & (\regs[0][5]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][5]~q ),
	.datad(\regs[1][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~560_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~560 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[5]~560 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \rfif.rdat2[5]~561 (
// Equation(s):
// \rfif.rdat2[5]~561_combout  = (Instr_IF_17 & ((\rfif.rdat2[5]~560_combout  & ((\regs[3][5]~q ))) # (!\rfif.rdat2[5]~560_combout  & (\regs[2][5]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[5]~560_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[2][5]~q ),
	.datac(\regs[3][5]~q ),
	.datad(\rfif.rdat2[5]~560_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~561_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~561 .lut_mask = 16'hF588;
defparam \rfif.rdat2[5]~561 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N25
dffeas \regs[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][5] .is_wysiwyg = "true";
defparam \regs[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N11
dffeas \regs[7][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][5] .is_wysiwyg = "true";
defparam \regs[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N27
dffeas \regs[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][5] .is_wysiwyg = "true";
defparam \regs[4][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N1
dffeas \regs[6][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][5] .is_wysiwyg = "true";
defparam \regs[6][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[5]~558 (
// Equation(s):
// \rfif.rdat2[5]~558_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[6][5]~q ))) # (!Instr_IF_17 & (\regs[4][5]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][5]~q ),
	.datad(\regs[6][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~558_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~558 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[5]~558 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[5]~559 (
// Equation(s):
// \rfif.rdat2[5]~559_combout  = (Instr_IF_16 & ((\rfif.rdat2[5]~558_combout  & ((\regs[7][5]~q ))) # (!\rfif.rdat2[5]~558_combout  & (\regs[5][5]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[5]~558_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][5]~q ),
	.datac(\regs[7][5]~q ),
	.datad(\rfif.rdat2[5]~558_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~559_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~559 .lut_mask = 16'hF588;
defparam \rfif.rdat2[5]~559 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[5]~562 (
// Equation(s):
// \rfif.rdat2[5]~562_combout  = (Instr_IF_18 & (((Instr_IF_19) # (\rfif.rdat2[5]~559_combout )))) # (!Instr_IF_18 & (\rfif.rdat2[5]~561_combout  & (!Instr_IF_19)))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[5]~561_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[5]~559_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~562_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~562 .lut_mask = 16'hAEA4;
defparam \rfif.rdat2[5]~562 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \rfif.rdat2[5]~565 (
// Equation(s):
// \rfif.rdat2[5]~565_combout  = (Instr_IF_19 & ((\rfif.rdat2[5]~562_combout  & ((\rfif.rdat2[5]~564_combout ))) # (!\rfif.rdat2[5]~562_combout  & (\rfif.rdat2[5]~557_combout )))) # (!Instr_IF_19 & (((\rfif.rdat2[5]~562_combout ))))

	.dataa(\rfif.rdat2[5]~557_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[5]~564_combout ),
	.datad(\rfif.rdat2[5]~562_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[5]~565_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[5]~565 .lut_mask = 16'hF388;
defparam \rfif.rdat2[5]~565 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N11
dffeas \regs[19][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][5] .is_wysiwyg = "true";
defparam \regs[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[5]~527 (
// Equation(s):
// \rfif.rdat1[5]~527_combout  = (Instr_IF_24 & ((Instr_IF_23) # ((\regs[27][5]~q )))) # (!Instr_IF_24 & (!Instr_IF_23 & ((\regs[19][5]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[27][5]~q ),
	.datad(\regs[19][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~527_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~527 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[5]~527 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \regs[23][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][5] .is_wysiwyg = "true";
defparam \regs[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[5]~528 (
// Equation(s):
// \rfif.rdat1[5]~528_combout  = (\rfif.rdat1[5]~527_combout  & ((\regs[31][5]~q ) # ((!Instr_IF_23)))) # (!\rfif.rdat1[5]~527_combout  & (((\regs[23][5]~q  & Instr_IF_23))))

	.dataa(\rfif.rdat1[5]~527_combout ),
	.datab(\regs[31][5]~q ),
	.datac(\regs[23][5]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~528_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~528 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[5]~528 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N27
dffeas \regs[29][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][5] .is_wysiwyg = "true";
defparam \regs[29][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas \regs[21][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][5] .is_wysiwyg = "true";
defparam \regs[21][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N13
dffeas \regs[25][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][5] .is_wysiwyg = "true";
defparam \regs[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[5]~520 (
// Equation(s):
// \rfif.rdat1[5]~520_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][5]~q ))) # (!Instr_IF_24 & (\regs[17][5]~q ))))

	.dataa(\regs[17][5]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[25][5]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~520_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~520 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[5]~520 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \rfif.rdat1[5]~521 (
// Equation(s):
// \rfif.rdat1[5]~521_combout  = (Instr_IF_23 & ((\rfif.rdat1[5]~520_combout  & (\regs[29][5]~q )) # (!\rfif.rdat1[5]~520_combout  & ((\regs[21][5]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[5]~520_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[29][5]~q ),
	.datac(\regs[21][5]~q ),
	.datad(\rfif.rdat1[5]~520_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~521_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~521 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[5]~521 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N13
dffeas \regs[26][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][5] .is_wysiwyg = "true";
defparam \regs[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[5]~523 (
// Equation(s):
// \rfif.rdat1[5]~523_combout  = (\rfif.rdat1[5]~522_combout  & (((\regs[30][5]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[5]~522_combout  & (Instr_IF_24 & ((\regs[26][5]~q ))))

	.dataa(\rfif.rdat1[5]~522_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[30][5]~q ),
	.datad(\regs[26][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~523_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~523 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[5]~523 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N8
cycloneive_lcell_comb \rfif.rdat1[5]~525 (
// Equation(s):
// \rfif.rdat1[5]~525_combout  = (\rfif.rdat1[5]~524_combout  & (((\regs[28][5]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[5]~524_combout  & (Instr_IF_24 & (\regs[24][5]~q )))

	.dataa(\rfif.rdat1[5]~524_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[24][5]~q ),
	.datad(\regs[28][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~525_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~525 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[5]~525 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N6
cycloneive_lcell_comb \rfif.rdat1[5]~526 (
// Equation(s):
// \rfif.rdat1[5]~526_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\rfif.rdat1[5]~523_combout )) # (!Instr_IF_22 & ((\rfif.rdat1[5]~525_combout )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\rfif.rdat1[5]~523_combout ),
	.datad(\rfif.rdat1[5]~525_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~526_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~526 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[5]~526 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[5]~530 (
// Equation(s):
// \rfif.rdat1[5]~530_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[5][5]~q ))) # (!Instr_IF_21 & (\regs[4][5]~q ))))

	.dataa(Instr_IF_22),
	.datab(\regs[4][5]~q ),
	.datac(\regs[5][5]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~530_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~530 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[5]~530 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \rfif.rdat1[5]~531 (
// Equation(s):
// \rfif.rdat1[5]~531_combout  = (Instr_IF_22 & ((\rfif.rdat1[5]~530_combout  & ((\regs[7][5]~q ))) # (!\rfif.rdat1[5]~530_combout  & (\regs[6][5]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[5]~530_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[5]~530_combout ),
	.datac(\regs[6][5]~q ),
	.datad(\regs[7][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~531_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~531 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[5]~531 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[5]~537 (
// Equation(s):
// \rfif.rdat1[5]~537_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[13][5]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & (\regs[12][5]~q )))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[12][5]~q ),
	.datad(\regs[13][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~537_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~537 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[5]~537 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \rfif.rdat1[5]~538 (
// Equation(s):
// \rfif.rdat1[5]~538_combout  = (Instr_IF_22 & ((\rfif.rdat1[5]~537_combout  & (\regs[15][5]~q )) # (!\rfif.rdat1[5]~537_combout  & ((\regs[14][5]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[5]~537_combout ))))

	.dataa(\regs[15][5]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[14][5]~q ),
	.datad(\rfif.rdat1[5]~537_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~538_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~538 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[5]~538 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[5]~534 (
// Equation(s):
// \rfif.rdat1[5]~534_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[2][5]~q ))) # (!Instr_IF_22 & (\regs[0][5]~q ))))

	.dataa(\regs[0][5]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[2][5]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~534_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~534 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[5]~534 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \rfif.rdat1[5]~535 (
// Equation(s):
// \rfif.rdat1[5]~535_combout  = (Instr_IF_21 & ((\rfif.rdat1[5]~534_combout  & (\regs[3][5]~q )) # (!\rfif.rdat1[5]~534_combout  & ((\regs[1][5]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[5]~534_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[3][5]~q ),
	.datac(\regs[1][5]~q ),
	.datad(\rfif.rdat1[5]~534_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~535_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~535 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[5]~535 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N4
cycloneive_lcell_comb \rfif.rdat1[5]~532 (
// Equation(s):
// \rfif.rdat1[5]~532_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][5]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\regs[8][5]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[10][5]~q ),
	.datad(\regs[8][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~532_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~532 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[5]~532 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N24
cycloneive_lcell_comb \rfif.rdat1[5]~533 (
// Equation(s):
// \rfif.rdat1[5]~533_combout  = (Instr_IF_21 & ((\rfif.rdat1[5]~532_combout  & ((\regs[11][5]~q ))) # (!\rfif.rdat1[5]~532_combout  & (\regs[9][5]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[5]~532_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[5]~532_combout ),
	.datac(\regs[9][5]~q ),
	.datad(\regs[11][5]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~533_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~533 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[5]~533 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N4
cycloneive_lcell_comb \rfif.rdat1[5]~536 (
// Equation(s):
// \rfif.rdat1[5]~536_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[5]~533_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[5]~535_combout ))))

	.dataa(\rfif.rdat1[5]~535_combout ),
	.datab(\rfif.rdat1[5]~533_combout ),
	.datac(Instr_IF_23),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[5]~536_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[5]~536 .lut_mask = 16'hFC0A;
defparam \rfif.rdat1[5]~536 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N15
dffeas \regs[0][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][4] .is_wysiwyg = "true";
defparam \regs[0][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N13
dffeas \regs[2][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][4] .is_wysiwyg = "true";
defparam \regs[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[4]~581 (
// Equation(s):
// \rfif.rdat2[4]~581_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[2][4]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[0][4]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[0][4]~q ),
	.datad(\regs[2][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~581_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~581 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[4]~581 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N15
dffeas \regs[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][4] .is_wysiwyg = "true";
defparam \regs[3][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N29
dffeas \regs[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][4] .is_wysiwyg = "true";
defparam \regs[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[4]~582 (
// Equation(s):
// \rfif.rdat2[4]~582_combout  = (Instr_IF_16 & ((\rfif.rdat2[4]~581_combout  & (\regs[3][4]~q )) # (!\rfif.rdat2[4]~581_combout  & ((\regs[1][4]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[4]~581_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[4]~581_combout ),
	.datac(\regs[3][4]~q ),
	.datad(\regs[1][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~582_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~582 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[4]~582 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[4]~583 (
// Equation(s):
// \rfif.rdat2[4]~583_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[4]~580_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[4]~582_combout )))))

	.dataa(\rfif.rdat2[4]~580_combout ),
	.datab(Instr_IF_18),
	.datac(\rfif.rdat2[4]~582_combout ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~583_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~583 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[4]~583 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N17
dffeas \regs[15][4] (
	.clk(!CLK),
	.d(input_a10),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][4] .is_wysiwyg = "true";
defparam \regs[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N31
dffeas \regs[14][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][4] .is_wysiwyg = "true";
defparam \regs[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N19
dffeas \regs[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][4] .is_wysiwyg = "true";
defparam \regs[13][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N5
dffeas \regs[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][4] .is_wysiwyg = "true";
defparam \regs[12][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N4
cycloneive_lcell_comb \rfif.rdat2[4]~584 (
// Equation(s):
// \rfif.rdat2[4]~584_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & (\regs[13][4]~q )) # (!Instr_IF_16 & ((\regs[12][4]~q )))))

	.dataa(Instr_IF_17),
	.datab(\regs[13][4]~q ),
	.datac(\regs[12][4]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~584_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~584 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[4]~584 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \rfif.rdat2[4]~585 (
// Equation(s):
// \rfif.rdat2[4]~585_combout  = (Instr_IF_17 & ((\rfif.rdat2[4]~584_combout  & (\regs[15][4]~q )) # (!\rfif.rdat2[4]~584_combout  & ((\regs[14][4]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[4]~584_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[15][4]~q ),
	.datac(\regs[14][4]~q ),
	.datad(\rfif.rdat2[4]~584_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~585_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~585 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[4]~585 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \regs[7][4]~feeder (
// Equation(s):
// \regs[7][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a10),
	.cin(gnd),
	.combout(\regs[7][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[7][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[7][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N15
dffeas \regs[7][4] (
	.clk(!CLK),
	.d(\regs[7][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][4] .is_wysiwyg = "true";
defparam \regs[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N27
dffeas \regs[6][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][4] .is_wysiwyg = "true";
defparam \regs[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N25
dffeas \regs[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][4] .is_wysiwyg = "true";
defparam \regs[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \regs[5][4]~feeder (
// Equation(s):
// \regs[5][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a10),
	.cin(gnd),
	.combout(\regs[5][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[5][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[5][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N11
dffeas \regs[5][4] (
	.clk(!CLK),
	.d(\regs[5][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][4] .is_wysiwyg = "true";
defparam \regs[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \rfif.rdat2[4]~577 (
// Equation(s):
// \rfif.rdat2[4]~577_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][4]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[4][4]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[4][4]~q ),
	.datad(\regs[5][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~577_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~577 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[4]~577 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \rfif.rdat2[4]~578 (
// Equation(s):
// \rfif.rdat2[4]~578_combout  = (Instr_IF_17 & ((\rfif.rdat2[4]~577_combout  & (\regs[7][4]~q )) # (!\rfif.rdat2[4]~577_combout  & ((\regs[6][4]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[4]~577_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[7][4]~q ),
	.datac(\regs[6][4]~q ),
	.datad(\rfif.rdat2[4]~577_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~578_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~578 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[4]~578 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[4]~586 (
// Equation(s):
// \rfif.rdat2[4]~586_combout  = (\rfif.rdat2[4]~583_combout  & ((\rfif.rdat2[4]~585_combout ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[4]~583_combout  & (((Instr_IF_18 & \rfif.rdat2[4]~578_combout ))))

	.dataa(\rfif.rdat2[4]~583_combout ),
	.datab(\rfif.rdat2[4]~585_combout ),
	.datac(Instr_IF_18),
	.datad(\rfif.rdat2[4]~578_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~586_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~586 .lut_mask = 16'hDA8A;
defparam \rfif.rdat2[4]~586 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N23
dffeas \regs[18][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][4] .is_wysiwyg = "true";
defparam \regs[18][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N21
dffeas \regs[22][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][4] .is_wysiwyg = "true";
defparam \regs[22][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \rfif.rdat2[4]~569 (
// Equation(s):
// \rfif.rdat2[4]~569_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][4]~q ))) # (!Instr_IF_18 & (\regs[18][4]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][4]~q ),
	.datad(\regs[22][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~569_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~569 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[4]~569 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N19
dffeas \regs[30][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][4] .is_wysiwyg = "true";
defparam \regs[30][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N13
dffeas \regs[26][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][4] .is_wysiwyg = "true";
defparam \regs[26][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[4]~570 (
// Equation(s):
// \rfif.rdat2[4]~570_combout  = (Instr_IF_19 & ((\rfif.rdat2[4]~569_combout  & (\regs[30][4]~q )) # (!\rfif.rdat2[4]~569_combout  & ((\regs[26][4]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[4]~569_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[4]~569_combout ),
	.datac(\regs[30][4]~q ),
	.datad(\regs[26][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~570_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~570 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[4]~570 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N21
dffeas \regs[24][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][4] .is_wysiwyg = "true";
defparam \regs[24][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N30
cycloneive_lcell_comb \regs[28][4]~feeder (
// Equation(s):
// \regs[28][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a10),
	.cin(gnd),
	.combout(\regs[28][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[28][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[28][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N31
dffeas \regs[28][4] (
	.clk(!CLK),
	.d(\regs[28][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][4] .is_wysiwyg = "true";
defparam \regs[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N19
dffeas \regs[16][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][4] .is_wysiwyg = "true";
defparam \regs[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[4]~571 (
// Equation(s):
// \rfif.rdat2[4]~571_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[20][4]~q )) # (!Instr_IF_18 & ((\regs[16][4]~q )))))

	.dataa(\regs[20][4]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[16][4]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~571_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~571 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[4]~571 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \rfif.rdat2[4]~572 (
// Equation(s):
// \rfif.rdat2[4]~572_combout  = (Instr_IF_19 & ((\rfif.rdat2[4]~571_combout  & ((\regs[28][4]~q ))) # (!\rfif.rdat2[4]~571_combout  & (\regs[24][4]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[4]~571_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[24][4]~q ),
	.datac(\regs[28][4]~q ),
	.datad(\rfif.rdat2[4]~571_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~572_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~572 .lut_mask = 16'hF588;
defparam \rfif.rdat2[4]~572 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \rfif.rdat2[4]~573 (
// Equation(s):
// \rfif.rdat2[4]~573_combout  = (Instr_IF_17 & ((\rfif.rdat2[4]~570_combout ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\rfif.rdat2[4]~572_combout  & !Instr_IF_16))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[4]~570_combout ),
	.datac(\rfif.rdat2[4]~572_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~573_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~573 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[4]~573 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \regs[21][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][4] .is_wysiwyg = "true";
defparam \regs[21][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N31
dffeas \regs[25][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][4] .is_wysiwyg = "true";
defparam \regs[25][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N31
dffeas \regs[17][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][4] .is_wysiwyg = "true";
defparam \regs[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \rfif.rdat2[4]~567 (
// Equation(s):
// \rfif.rdat2[4]~567_combout  = (Instr_IF_19 & ((Instr_IF_18) # ((\regs[25][4]~q )))) # (!Instr_IF_19 & (!Instr_IF_18 & ((\regs[17][4]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[25][4]~q ),
	.datad(\regs[17][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~567_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~567 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[4]~567 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \rfif.rdat2[4]~568 (
// Equation(s):
// \rfif.rdat2[4]~568_combout  = (Instr_IF_18 & ((\rfif.rdat2[4]~567_combout  & (\regs[29][4]~q )) # (!\rfif.rdat2[4]~567_combout  & ((\regs[21][4]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[4]~567_combout ))))

	.dataa(\regs[29][4]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[21][4]~q ),
	.datad(\rfif.rdat2[4]~567_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~568_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~568 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[4]~568 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N13
dffeas \regs[23][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][4] .is_wysiwyg = "true";
defparam \regs[23][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \regs[31][4]~feeder (
// Equation(s):
// \regs[31][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a10),
	.cin(gnd),
	.combout(\regs[31][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[31][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[31][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N17
dffeas \regs[31][4] (
	.clk(!CLK),
	.d(\regs[31][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][4] .is_wysiwyg = "true";
defparam \regs[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[4]~575 (
// Equation(s):
// \rfif.rdat2[4]~575_combout  = (\rfif.rdat2[4]~574_combout  & (((\regs[31][4]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[4]~574_combout  & (\regs[23][4]~q  & (Instr_IF_18)))

	.dataa(\rfif.rdat2[4]~574_combout ),
	.datab(\regs[23][4]~q ),
	.datac(Instr_IF_18),
	.datad(\regs[31][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~575_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~575 .lut_mask = 16'hEA4A;
defparam \rfif.rdat2[4]~575 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[4]~576 (
// Equation(s):
// \rfif.rdat2[4]~576_combout  = (\rfif.rdat2[4]~573_combout  & (((\rfif.rdat2[4]~575_combout )) # (!Instr_IF_16))) # (!\rfif.rdat2[4]~573_combout  & (Instr_IF_16 & (\rfif.rdat2[4]~568_combout )))

	.dataa(\rfif.rdat2[4]~573_combout ),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[4]~568_combout ),
	.datad(\rfif.rdat2[4]~575_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[4]~576_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[4]~576 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[4]~576 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N20
cycloneive_lcell_comb \regs[20][4]~feeder (
// Equation(s):
// \regs[20][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a10),
	.cin(gnd),
	.combout(\regs[20][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[20][4]~feeder .lut_mask = 16'hFF00;
defparam \regs[20][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N21
dffeas \regs[20][4] (
	.clk(!CLK),
	.d(\regs[20][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][4] .is_wysiwyg = "true";
defparam \regs[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[4]~544 (
// Equation(s):
// \rfif.rdat1[4]~544_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][4]~q ))) # (!Instr_IF_24 & (\regs[16][4]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][4]~q ),
	.datac(\regs[24][4]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~544_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~544 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[4]~544 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \rfif.rdat1[4]~545 (
// Equation(s):
// \rfif.rdat1[4]~545_combout  = (Instr_IF_23 & ((\rfif.rdat1[4]~544_combout  & ((\regs[28][4]~q ))) # (!\rfif.rdat1[4]~544_combout  & (\regs[20][4]~q )))) # (!Instr_IF_23 & (((\rfif.rdat1[4]~544_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[20][4]~q ),
	.datac(\regs[28][4]~q ),
	.datad(\rfif.rdat1[4]~544_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~545_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~545 .lut_mask = 16'hF588;
defparam \rfif.rdat1[4]~545 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \rfif.rdat1[4]~542 (
// Equation(s):
// \rfif.rdat1[4]~542_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[21][4]~q ))) # (!Instr_IF_23 & (\regs[17][4]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[17][4]~q ),
	.datad(\regs[21][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~542_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~542 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[4]~542 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N1
dffeas \regs[29][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][4] .is_wysiwyg = "true";
defparam \regs[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[4]~543 (
// Equation(s):
// \rfif.rdat1[4]~543_combout  = (\rfif.rdat1[4]~542_combout  & (((\regs[29][4]~q ) # (!Instr_IF_24)))) # (!\rfif.rdat1[4]~542_combout  & (\regs[25][4]~q  & ((Instr_IF_24))))

	.dataa(\regs[25][4]~q ),
	.datab(\rfif.rdat1[4]~542_combout ),
	.datac(\regs[29][4]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~543_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~543 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[4]~543 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \rfif.rdat1[4]~546 (
// Equation(s):
// \rfif.rdat1[4]~546_combout  = (Instr_IF_21 & (((Instr_IF_22) # (\rfif.rdat1[4]~543_combout )))) # (!Instr_IF_21 & (\rfif.rdat1[4]~545_combout  & (!Instr_IF_22)))

	.dataa(\rfif.rdat1[4]~545_combout ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[4]~543_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~546_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~546 .lut_mask = 16'hCEC2;
defparam \rfif.rdat1[4]~546 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N19
dffeas \regs[27][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][4] .is_wysiwyg = "true";
defparam \regs[27][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[4]~547 (
// Equation(s):
// \rfif.rdat1[4]~547_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][4]~q ))) # (!Instr_IF_23 & (\regs[19][4]~q ))))

	.dataa(\regs[19][4]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[23][4]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~547_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~547 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[4]~547 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \rfif.rdat1[4]~548 (
// Equation(s):
// \rfif.rdat1[4]~548_combout  = (Instr_IF_24 & ((\rfif.rdat1[4]~547_combout  & (\regs[31][4]~q )) # (!\rfif.rdat1[4]~547_combout  & ((\regs[27][4]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[4]~547_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[31][4]~q ),
	.datac(\regs[27][4]~q ),
	.datad(\rfif.rdat1[4]~547_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~548_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~548 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[4]~548 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[4]~540 (
// Equation(s):
// \rfif.rdat1[4]~540_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][4]~q )) # (!Instr_IF_24 & ((\regs[18][4]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][4]~q ),
	.datad(\regs[18][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~540_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~540 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[4]~540 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[4]~541 (
// Equation(s):
// \rfif.rdat1[4]~541_combout  = (Instr_IF_23 & ((\rfif.rdat1[4]~540_combout  & (\regs[30][4]~q )) # (!\rfif.rdat1[4]~540_combout  & ((\regs[22][4]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[4]~540_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[30][4]~q ),
	.datac(\regs[22][4]~q ),
	.datad(\rfif.rdat1[4]~540_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~541_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~541 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[4]~541 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[4]~554 (
// Equation(s):
// \rfif.rdat1[4]~554_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][4]~q )) # (!Instr_IF_21 & ((\regs[0][4]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][4]~q ),
	.datad(\regs[0][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~554_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~554 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[4]~554 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \rfif.rdat1[4]~555 (
// Equation(s):
// \rfif.rdat1[4]~555_combout  = (Instr_IF_22 & ((\rfif.rdat1[4]~554_combout  & ((\regs[3][4]~q ))) # (!\rfif.rdat1[4]~554_combout  & (\regs[2][4]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[4]~554_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[4]~554_combout ),
	.datac(\regs[2][4]~q ),
	.datad(\regs[3][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~555_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~555 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[4]~555 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \rfif.rdat1[4]~552 (
// Equation(s):
// \rfif.rdat1[4]~552_combout  = (Instr_IF_22 & ((\regs[6][4]~q ) # ((Instr_IF_21)))) # (!Instr_IF_22 & (((\regs[4][4]~q  & !Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[6][4]~q ),
	.datac(\regs[4][4]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~552_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~552 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[4]~552 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \rfif.rdat1[4]~553 (
// Equation(s):
// \rfif.rdat1[4]~553_combout  = (Instr_IF_21 & ((\rfif.rdat1[4]~552_combout  & (\regs[7][4]~q )) # (!\rfif.rdat1[4]~552_combout  & ((\regs[5][4]~q ))))) # (!Instr_IF_21 & (\rfif.rdat1[4]~552_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[4]~552_combout ),
	.datac(\regs[7][4]~q ),
	.datad(\regs[5][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~553_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~553 .lut_mask = 16'hE6C4;
defparam \rfif.rdat1[4]~553 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N12
cycloneive_lcell_comb \rfif.rdat1[4]~556 (
// Equation(s):
// \rfif.rdat1[4]~556_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\rfif.rdat1[4]~553_combout )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\rfif.rdat1[4]~555_combout )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[4]~555_combout ),
	.datad(\rfif.rdat1[4]~553_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~556_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~556 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[4]~556 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \rfif.rdat1[4]~557 (
// Equation(s):
// \rfif.rdat1[4]~557_combout  = (Instr_IF_22 & (((\regs[14][4]~q ) # (Instr_IF_21)))) # (!Instr_IF_22 & (\regs[12][4]~q  & ((!Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[12][4]~q ),
	.datac(\regs[14][4]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~557_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~557 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[4]~557 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N18
cycloneive_lcell_comb \rfif.rdat1[4]~558 (
// Equation(s):
// \rfif.rdat1[4]~558_combout  = (\rfif.rdat1[4]~557_combout  & (((\regs[15][4]~q )) # (!Instr_IF_21))) # (!\rfif.rdat1[4]~557_combout  & (Instr_IF_21 & (\regs[13][4]~q )))

	.dataa(\rfif.rdat1[4]~557_combout ),
	.datab(Instr_IF_21),
	.datac(\regs[13][4]~q ),
	.datad(\regs[15][4]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~558_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~558 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[4]~558 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N14
cycloneive_lcell_comb \regs[11][4]~feeder (
// Equation(s):
// \regs[11][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[11][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[11][4]~feeder .lut_mask = 16'hF0F0;
defparam \regs[11][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N15
dffeas \regs[11][4] (
	.clk(!CLK),
	.d(\regs[11][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][4] .is_wysiwyg = "true";
defparam \regs[11][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N24
cycloneive_lcell_comb \regs[10][4]~feeder (
// Equation(s):
// \regs[10][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[10][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[10][4]~feeder .lut_mask = 16'hF0F0;
defparam \regs[10][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N25
dffeas \regs[10][4] (
	.clk(!CLK),
	.d(\regs[10][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][4] .is_wysiwyg = "true";
defparam \regs[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N4
cycloneive_lcell_comb \regs[9][4]~feeder (
// Equation(s):
// \regs[9][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[9][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[9][4]~feeder .lut_mask = 16'hF0F0;
defparam \regs[9][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N5
dffeas \regs[9][4] (
	.clk(!CLK),
	.d(\regs[9][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][4] .is_wysiwyg = "true";
defparam \regs[9][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N6
cycloneive_lcell_comb \regs[8][4]~feeder (
// Equation(s):
// \regs[8][4]~feeder_combout  = \input_a~123_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a10),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[8][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[8][4]~feeder .lut_mask = 16'hF0F0;
defparam \regs[8][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N7
dffeas \regs[8][4] (
	.clk(!CLK),
	.d(\regs[8][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][4] .is_wysiwyg = "true";
defparam \regs[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N0
cycloneive_lcell_comb \rfif.rdat1[4]~550 (
// Equation(s):
// \rfif.rdat1[4]~550_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[9][4]~q )) # (!Instr_IF_21 & ((\regs[8][4]~q )))))

	.dataa(Instr_IF_22),
	.datab(\regs[9][4]~q ),
	.datac(\regs[8][4]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~550_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~550 .lut_mask = 16'hEE50;
defparam \rfif.rdat1[4]~550 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N2
cycloneive_lcell_comb \rfif.rdat1[4]~551 (
// Equation(s):
// \rfif.rdat1[4]~551_combout  = (Instr_IF_22 & ((\rfif.rdat1[4]~550_combout  & (\regs[11][4]~q )) # (!\rfif.rdat1[4]~550_combout  & ((\regs[10][4]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[4]~550_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[11][4]~q ),
	.datac(\regs[10][4]~q ),
	.datad(\rfif.rdat1[4]~550_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[4]~551_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[4]~551 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[4]~551 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N17
dffeas \regs[22][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][3] .is_wysiwyg = "true";
defparam \regs[22][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N31
dffeas \regs[18][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][3] .is_wysiwyg = "true";
defparam \regs[18][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N29
dffeas \regs[26][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][3] .is_wysiwyg = "true";
defparam \regs[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \rfif.rdat2[3]~588 (
// Equation(s):
// \rfif.rdat2[3]~588_combout  = (Instr_IF_19 & (((\regs[26][3]~q ) # (Instr_IF_18)))) # (!Instr_IF_19 & (\regs[18][3]~q  & ((!Instr_IF_18))))

	.dataa(Instr_IF_19),
	.datab(\regs[18][3]~q ),
	.datac(\regs[26][3]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~588_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~588 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[3]~588 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \rfif.rdat2[3]~589 (
// Equation(s):
// \rfif.rdat2[3]~589_combout  = (Instr_IF_18 & ((\rfif.rdat2[3]~588_combout  & (\regs[30][3]~q )) # (!\rfif.rdat2[3]~588_combout  & ((\regs[22][3]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[3]~588_combout ))))

	.dataa(\regs[30][3]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[22][3]~q ),
	.datad(\rfif.rdat2[3]~588_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~589_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~589 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[3]~589 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \regs[31][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][3] .is_wysiwyg = "true";
defparam \regs[31][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N25
dffeas \regs[27][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][3] .is_wysiwyg = "true";
defparam \regs[27][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \rfif.rdat2[3]~596 (
// Equation(s):
// \rfif.rdat2[3]~596_combout  = (\rfif.rdat2[3]~595_combout  & (((\regs[31][3]~q )) # (!Instr_IF_19))) # (!\rfif.rdat2[3]~595_combout  & (Instr_IF_19 & ((\regs[27][3]~q ))))

	.dataa(\rfif.rdat2[3]~595_combout ),
	.datab(Instr_IF_19),
	.datac(\regs[31][3]~q ),
	.datad(\regs[27][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~596_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~596 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[3]~596 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N17
dffeas \regs[25][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][3] .is_wysiwyg = "true";
defparam \regs[25][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N23
dffeas \regs[29][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][3] .is_wysiwyg = "true";
defparam \regs[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N27
dffeas \regs[17][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][3] .is_wysiwyg = "true";
defparam \regs[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \rfif.rdat2[3]~590 (
// Equation(s):
// \rfif.rdat2[3]~590_combout  = (Instr_IF_19 & (((Instr_IF_18)))) # (!Instr_IF_19 & ((Instr_IF_18 & (\regs[21][3]~q )) # (!Instr_IF_18 & ((\regs[17][3]~q )))))

	.dataa(\regs[21][3]~q ),
	.datab(Instr_IF_19),
	.datac(\regs[17][3]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~590_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~590 .lut_mask = 16'hEE30;
defparam \rfif.rdat2[3]~590 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \rfif.rdat2[3]~591 (
// Equation(s):
// \rfif.rdat2[3]~591_combout  = (Instr_IF_19 & ((\rfif.rdat2[3]~590_combout  & ((\regs[29][3]~q ))) # (!\rfif.rdat2[3]~590_combout  & (\regs[25][3]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[3]~590_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[25][3]~q ),
	.datac(\regs[29][3]~q ),
	.datad(\rfif.rdat2[3]~590_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~591_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~591 .lut_mask = 16'hF588;
defparam \rfif.rdat2[3]~591 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N19
dffeas \regs[28][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][3] .is_wysiwyg = "true";
defparam \regs[28][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N3
dffeas \regs[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][3] .is_wysiwyg = "true";
defparam \regs[16][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N29
dffeas \regs[24][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][3] .is_wysiwyg = "true";
defparam \regs[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[3]~592 (
// Equation(s):
// \rfif.rdat2[3]~592_combout  = (Instr_IF_18 & (Instr_IF_19)) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[24][3]~q ))) # (!Instr_IF_19 & (\regs[16][3]~q ))))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][3]~q ),
	.datad(\regs[24][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~592_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~592 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[3]~592 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N18
cycloneive_lcell_comb \rfif.rdat2[3]~593 (
// Equation(s):
// \rfif.rdat2[3]~593_combout  = (Instr_IF_18 & ((\rfif.rdat2[3]~592_combout  & ((\regs[28][3]~q ))) # (!\rfif.rdat2[3]~592_combout  & (\regs[20][3]~q )))) # (!Instr_IF_18 & (((\rfif.rdat2[3]~592_combout ))))

	.dataa(\regs[20][3]~q ),
	.datab(Instr_IF_18),
	.datac(\regs[28][3]~q ),
	.datad(\rfif.rdat2[3]~592_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~593_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~593 .lut_mask = 16'hF388;
defparam \rfif.rdat2[3]~593 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[3]~594 (
// Equation(s):
// \rfif.rdat2[3]~594_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & (\rfif.rdat2[3]~591_combout )) # (!Instr_IF_16 & ((\rfif.rdat2[3]~593_combout )))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[3]~591_combout ),
	.datad(\rfif.rdat2[3]~593_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~594_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~594 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[3]~594 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[3]~597 (
// Equation(s):
// \rfif.rdat2[3]~597_combout  = (\rfif.rdat2[3]~594_combout  & (((\rfif.rdat2[3]~596_combout ) # (!Instr_IF_17)))) # (!\rfif.rdat2[3]~594_combout  & (\rfif.rdat2[3]~589_combout  & ((Instr_IF_17))))

	.dataa(\rfif.rdat2[3]~589_combout ),
	.datab(\rfif.rdat2[3]~596_combout ),
	.datac(\rfif.rdat2[3]~594_combout ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~597_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~597 .lut_mask = 16'hCAF0;
defparam \rfif.rdat2[3]~597 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N29
dffeas \regs[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][3] .is_wysiwyg = "true";
defparam \regs[2][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N3
dffeas \regs[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][3] .is_wysiwyg = "true";
defparam \regs[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \rfif.rdat2[3]~603 (
// Equation(s):
// \rfif.rdat2[3]~603_combout  = (\rfif.rdat2[3]~602_combout  & (((\regs[3][3]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[3]~602_combout  & (\regs[2][3]~q  & ((Instr_IF_17))))

	.dataa(\rfif.rdat2[3]~602_combout ),
	.datab(\regs[2][3]~q ),
	.datac(\regs[3][3]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~603_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~603 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[3]~603 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[3]~604 (
// Equation(s):
// \rfif.rdat2[3]~604_combout  = (Instr_IF_18 & ((\rfif.rdat2[3]~601_combout ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((!Instr_IF_19 & \rfif.rdat2[3]~603_combout ))))

	.dataa(\rfif.rdat2[3]~601_combout ),
	.datab(Instr_IF_18),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[3]~603_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~604_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~604 .lut_mask = 16'hCBC8;
defparam \rfif.rdat2[3]~604 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N11
dffeas \regs[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][3] .is_wysiwyg = "true";
defparam \regs[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N19
dffeas \regs[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][3] .is_wysiwyg = "true";
defparam \regs[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N18
cycloneive_lcell_comb \rfif.rdat2[3]~605 (
// Equation(s):
// \rfif.rdat2[3]~605_combout  = (Instr_IF_17 & ((\regs[14][3]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\regs[12][3]~q  & !Instr_IF_16))))

	.dataa(Instr_IF_17),
	.datab(\regs[14][3]~q ),
	.datac(\regs[12][3]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~605_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~605 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[3]~605 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N29
dffeas \regs[15][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][3] .is_wysiwyg = "true";
defparam \regs[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N28
cycloneive_lcell_comb \rfif.rdat2[3]~606 (
// Equation(s):
// \rfif.rdat2[3]~606_combout  = (\rfif.rdat2[3]~605_combout  & (((\regs[15][3]~q ) # (!Instr_IF_16)))) # (!\rfif.rdat2[3]~605_combout  & (\regs[13][3]~q  & ((Instr_IF_16))))

	.dataa(\regs[13][3]~q ),
	.datab(\rfif.rdat2[3]~605_combout ),
	.datac(\regs[15][3]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~606_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~606 .lut_mask = 16'hE2CC;
defparam \rfif.rdat2[3]~606 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N9
dffeas \regs[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][3] .is_wysiwyg = "true";
defparam \regs[10][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N19
dffeas \regs[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][3] .is_wysiwyg = "true";
defparam \regs[11][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N8
cycloneive_lcell_comb \rfif.rdat2[3]~599 (
// Equation(s):
// \rfif.rdat2[3]~599_combout  = (\rfif.rdat2[3]~598_combout  & (((\regs[11][3]~q )) # (!Instr_IF_17))) # (!\rfif.rdat2[3]~598_combout  & (Instr_IF_17 & (\regs[10][3]~q )))

	.dataa(\rfif.rdat2[3]~598_combout ),
	.datab(Instr_IF_17),
	.datac(\regs[10][3]~q ),
	.datad(\regs[11][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~599_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~599 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[3]~599 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \rfif.rdat2[3]~607 (
// Equation(s):
// \rfif.rdat2[3]~607_combout  = (\rfif.rdat2[3]~604_combout  & (((\rfif.rdat2[3]~606_combout )) # (!Instr_IF_19))) # (!\rfif.rdat2[3]~604_combout  & (Instr_IF_19 & ((\rfif.rdat2[3]~599_combout ))))

	.dataa(\rfif.rdat2[3]~604_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[3]~606_combout ),
	.datad(\rfif.rdat2[3]~599_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[3]~607_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[3]~607 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[3]~607 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \regs[23][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][3] .is_wysiwyg = "true";
defparam \regs[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \regs[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][3] .is_wysiwyg = "true";
defparam \regs[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[3]~567 (
// Equation(s):
// \rfif.rdat1[3]~567_combout  = (Instr_IF_24 & (((\regs[27][3]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[19][3]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[19][3]~q ),
	.datac(\regs[27][3]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~567_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~567 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[3]~567 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[3]~568 (
// Equation(s):
// \rfif.rdat1[3]~568_combout  = (Instr_IF_23 & ((\rfif.rdat1[3]~567_combout  & (\regs[31][3]~q )) # (!\rfif.rdat1[3]~567_combout  & ((\regs[23][3]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[3]~567_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[31][3]~q ),
	.datac(\regs[23][3]~q ),
	.datad(\rfif.rdat1[3]~567_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~568_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~568 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[3]~568 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \rfif.rdat1[3]~560 (
// Equation(s):
// \rfif.rdat1[3]~560_combout  = (Instr_IF_24 & (((\regs[25][3]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[17][3]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[17][3]~q ),
	.datac(\regs[25][3]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~560_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~560 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[3]~560 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N13
dffeas \regs[21][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][3] .is_wysiwyg = "true";
defparam \regs[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N12
cycloneive_lcell_comb \rfif.rdat1[3]~561 (
// Equation(s):
// \rfif.rdat1[3]~561_combout  = (\rfif.rdat1[3]~560_combout  & (((\regs[29][3]~q )) # (!Instr_IF_23))) # (!\rfif.rdat1[3]~560_combout  & (Instr_IF_23 & (\regs[21][3]~q )))

	.dataa(\rfif.rdat1[3]~560_combout ),
	.datab(Instr_IF_23),
	.datac(\regs[21][3]~q ),
	.datad(\regs[29][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~561_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~561 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[3]~561 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N11
dffeas \regs[30][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][3] .is_wysiwyg = "true";
defparam \regs[30][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \rfif.rdat1[3]~563 (
// Equation(s):
// \rfif.rdat1[3]~563_combout  = (\rfif.rdat1[3]~562_combout  & (((\regs[30][3]~q )) # (!Instr_IF_24))) # (!\rfif.rdat1[3]~562_combout  & (Instr_IF_24 & ((\regs[26][3]~q ))))

	.dataa(\rfif.rdat1[3]~562_combout ),
	.datab(Instr_IF_24),
	.datac(\regs[30][3]~q ),
	.datad(\regs[26][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~563_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~563 .lut_mask = 16'hE6A2;
defparam \rfif.rdat1[3]~563 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[3]~565 (
// Equation(s):
// \rfif.rdat1[3]~565_combout  = (\rfif.rdat1[3]~564_combout  & ((\regs[28][3]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[3]~564_combout  & (((\regs[24][3]~q  & Instr_IF_24))))

	.dataa(\rfif.rdat1[3]~564_combout ),
	.datab(\regs[28][3]~q ),
	.datac(\regs[24][3]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~565_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~565 .lut_mask = 16'hD8AA;
defparam \rfif.rdat1[3]~565 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \rfif.rdat1[3]~566 (
// Equation(s):
// \rfif.rdat1[3]~566_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\rfif.rdat1[3]~563_combout )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\rfif.rdat1[3]~565_combout ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[3]~563_combout ),
	.datad(\rfif.rdat1[3]~565_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~566_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~566 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[3]~566 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N21
dffeas \regs[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][3] .is_wysiwyg = "true";
defparam \regs[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[3]~570 (
// Equation(s):
// \rfif.rdat1[3]~570_combout  = (Instr_IF_21 & (((\regs[5][3]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[4][3]~q  & ((!Instr_IF_22))))

	.dataa(\regs[4][3]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][3]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~570_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~570 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[3]~570 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N21
dffeas \regs[6][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][3] .is_wysiwyg = "true";
defparam \regs[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N3
dffeas \regs[7][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][3] .is_wysiwyg = "true";
defparam \regs[7][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[3]~571 (
// Equation(s):
// \rfif.rdat1[3]~571_combout  = (Instr_IF_22 & ((\rfif.rdat1[3]~570_combout  & ((\regs[7][3]~q ))) # (!\rfif.rdat1[3]~570_combout  & (\regs[6][3]~q )))) # (!Instr_IF_22 & (\rfif.rdat1[3]~570_combout ))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[3]~570_combout ),
	.datac(\regs[6][3]~q ),
	.datad(\regs[7][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~571_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~571 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[3]~571 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[3]~574 (
// Equation(s):
// \rfif.rdat1[3]~574_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[2][3]~q ))) # (!Instr_IF_22 & (\regs[0][3]~q ))))

	.dataa(\regs[0][3]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[2][3]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~574_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~574 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[3]~574 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N1
dffeas \regs[1][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][3] .is_wysiwyg = "true";
defparam \regs[1][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N0
cycloneive_lcell_comb \rfif.rdat1[3]~575 (
// Equation(s):
// \rfif.rdat1[3]~575_combout  = (Instr_IF_21 & ((\rfif.rdat1[3]~574_combout  & ((\regs[3][3]~q ))) # (!\rfif.rdat1[3]~574_combout  & (\regs[1][3]~q )))) # (!Instr_IF_21 & (\rfif.rdat1[3]~574_combout ))

	.dataa(Instr_IF_21),
	.datab(\rfif.rdat1[3]~574_combout ),
	.datac(\regs[1][3]~q ),
	.datad(\regs[3][3]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~575_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~575 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[3]~575 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N25
dffeas \regs[9][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][3] .is_wysiwyg = "true";
defparam \regs[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N3
dffeas \regs[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][3] .is_wysiwyg = "true";
defparam \regs[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N2
cycloneive_lcell_comb \rfif.rdat1[3]~572 (
// Equation(s):
// \rfif.rdat1[3]~572_combout  = (Instr_IF_22 & ((\regs[10][3]~q ) # ((Instr_IF_21)))) # (!Instr_IF_22 & (((\regs[8][3]~q  & !Instr_IF_21))))

	.dataa(Instr_IF_22),
	.datab(\regs[10][3]~q ),
	.datac(\regs[8][3]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~572_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~572 .lut_mask = 16'hAAD8;
defparam \rfif.rdat1[3]~572 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N18
cycloneive_lcell_comb \rfif.rdat1[3]~573 (
// Equation(s):
// \rfif.rdat1[3]~573_combout  = (Instr_IF_21 & ((\rfif.rdat1[3]~572_combout  & ((\regs[11][3]~q ))) # (!\rfif.rdat1[3]~572_combout  & (\regs[9][3]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[3]~572_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[9][3]~q ),
	.datac(\regs[11][3]~q ),
	.datad(\rfif.rdat1[3]~572_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~573_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~573 .lut_mask = 16'hF588;
defparam \rfif.rdat1[3]~573 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \rfif.rdat1[3]~576 (
// Equation(s):
// \rfif.rdat1[3]~576_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\rfif.rdat1[3]~573_combout ))) # (!Instr_IF_24 & (\rfif.rdat1[3]~575_combout ))))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[3]~575_combout ),
	.datac(Instr_IF_24),
	.datad(\rfif.rdat1[3]~573_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~576_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~576 .lut_mask = 16'hF4A4;
defparam \rfif.rdat1[3]~576 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N5
dffeas \regs[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][3] .is_wysiwyg = "true";
defparam \regs[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[3]~577 (
// Equation(s):
// \rfif.rdat1[3]~577_combout  = (Instr_IF_21 & (((\regs[13][3]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[12][3]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[12][3]~q ),
	.datac(\regs[13][3]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~577_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~577 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[3]~577 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \rfif.rdat1[3]~578 (
// Equation(s):
// \rfif.rdat1[3]~578_combout  = (\rfif.rdat1[3]~577_combout  & ((\regs[15][3]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[3]~577_combout  & (((\regs[14][3]~q  & Instr_IF_22))))

	.dataa(\regs[15][3]~q ),
	.datab(\rfif.rdat1[3]~577_combout ),
	.datac(\regs[14][3]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[3]~578_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[3]~578 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[3]~578 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N23
dffeas \regs[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][2] .is_wysiwyg = "true";
defparam \regs[5][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N3
dffeas \regs[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][2] .is_wysiwyg = "true";
defparam \regs[4][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \rfif.rdat2[2]~619 (
// Equation(s):
// \rfif.rdat2[2]~619_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[5][2]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & ((\regs[4][2]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[5][2]~q ),
	.datad(\regs[4][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~619_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~619 .lut_mask = 16'hB9A8;
defparam \rfif.rdat2[2]~619 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N29
dffeas \regs[6][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][2] .is_wysiwyg = "true";
defparam \regs[6][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \rfif.rdat2[2]~620 (
// Equation(s):
// \rfif.rdat2[2]~620_combout  = (\rfif.rdat2[2]~619_combout  & ((\regs[7][2]~q ) # ((!Instr_IF_17)))) # (!\rfif.rdat2[2]~619_combout  & (((\regs[6][2]~q  & Instr_IF_17))))

	.dataa(\regs[7][2]~q ),
	.datab(\rfif.rdat2[2]~619_combout ),
	.datac(\regs[6][2]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~620_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~620 .lut_mask = 16'hB8CC;
defparam \rfif.rdat2[2]~620 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N11
dffeas \regs[8][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][2] .is_wysiwyg = "true";
defparam \regs[8][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N13
dffeas \regs[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][2] .is_wysiwyg = "true";
defparam \regs[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \rfif.rdat2[2]~621 (
// Equation(s):
// \rfif.rdat2[2]~621_combout  = (Instr_IF_17 & ((Instr_IF_16) # ((\regs[10][2]~q )))) # (!Instr_IF_17 & (!Instr_IF_16 & (\regs[8][2]~q )))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[8][2]~q ),
	.datad(\regs[10][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~621_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~621 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[2]~621 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N27
dffeas \regs[11][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][2] .is_wysiwyg = "true";
defparam \regs[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N21
dffeas \regs[9][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][2] .is_wysiwyg = "true";
defparam \regs[9][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \rfif.rdat2[2]~622 (
// Equation(s):
// \rfif.rdat2[2]~622_combout  = (Instr_IF_16 & ((\rfif.rdat2[2]~621_combout  & (\regs[11][2]~q )) # (!\rfif.rdat2[2]~621_combout  & ((\regs[9][2]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[2]~621_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[2]~621_combout ),
	.datac(\regs[11][2]~q ),
	.datad(\regs[9][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~622_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~622 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[2]~622 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N15
dffeas \regs[2][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][2] .is_wysiwyg = "true";
defparam \regs[2][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N17
dffeas \regs[0][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][2] .is_wysiwyg = "true";
defparam \regs[0][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \rfif.rdat2[2]~623 (
// Equation(s):
// \rfif.rdat2[2]~623_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[2][2]~q )) # (!Instr_IF_17 & ((\regs[0][2]~q )))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[2][2]~q ),
	.datad(\regs[0][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~623_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~623 .lut_mask = 16'hD9C8;
defparam \rfif.rdat2[2]~623 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N23
dffeas \regs[3][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][2] .is_wysiwyg = "true";
defparam \regs[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \regs[1][2]~feeder (
// Equation(s):
// \regs[1][2]~feeder_combout  = \input_a~129_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a12),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[1][2]~feeder .lut_mask = 16'hF0F0;
defparam \regs[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N21
dffeas \regs[1][2] (
	.clk(!CLK),
	.d(\regs[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][2] .is_wysiwyg = "true";
defparam \regs[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \rfif.rdat2[2]~624 (
// Equation(s):
// \rfif.rdat2[2]~624_combout  = (Instr_IF_16 & ((\rfif.rdat2[2]~623_combout  & (\regs[3][2]~q )) # (!\rfif.rdat2[2]~623_combout  & ((\regs[1][2]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[2]~623_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[2]~623_combout ),
	.datac(\regs[3][2]~q ),
	.datad(\regs[1][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~624_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~624 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[2]~624 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \rfif.rdat2[2]~625 (
// Equation(s):
// \rfif.rdat2[2]~625_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & (\rfif.rdat2[2]~622_combout )) # (!Instr_IF_19 & ((\rfif.rdat2[2]~624_combout )))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[2]~622_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[2]~624_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~625_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~625 .lut_mask = 16'hE5E0;
defparam \rfif.rdat2[2]~625 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N3
dffeas \regs[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][2] .is_wysiwyg = "true";
defparam \regs[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N7
dffeas \regs[13][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][2] .is_wysiwyg = "true";
defparam \regs[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N2
cycloneive_lcell_comb \rfif.rdat2[2]~626 (
// Equation(s):
// \rfif.rdat2[2]~626_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[13][2]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[12][2]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[12][2]~q ),
	.datad(\regs[13][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~626_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~626 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[2]~626 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N17
dffeas \regs[15][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][2] .is_wysiwyg = "true";
defparam \regs[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N13
dffeas \regs[14][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][2] .is_wysiwyg = "true";
defparam \regs[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N16
cycloneive_lcell_comb \rfif.rdat2[2]~627 (
// Equation(s):
// \rfif.rdat2[2]~627_combout  = (Instr_IF_17 & ((\rfif.rdat2[2]~626_combout  & (\regs[15][2]~q )) # (!\rfif.rdat2[2]~626_combout  & ((\regs[14][2]~q ))))) # (!Instr_IF_17 & (\rfif.rdat2[2]~626_combout ))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[2]~626_combout ),
	.datac(\regs[15][2]~q ),
	.datad(\regs[14][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~627_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~627 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[2]~627 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[2]~628 (
// Equation(s):
// \rfif.rdat2[2]~628_combout  = (Instr_IF_18 & ((\rfif.rdat2[2]~625_combout  & ((\rfif.rdat2[2]~627_combout ))) # (!\rfif.rdat2[2]~625_combout  & (\rfif.rdat2[2]~620_combout )))) # (!Instr_IF_18 & (((\rfif.rdat2[2]~625_combout ))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[2]~620_combout ),
	.datac(\rfif.rdat2[2]~625_combout ),
	.datad(\rfif.rdat2[2]~627_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~628_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~628 .lut_mask = 16'hF858;
defparam \rfif.rdat2[2]~628 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N9
dffeas \regs[23][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][2] .is_wysiwyg = "true";
defparam \regs[23][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N13
dffeas \regs[31][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][2] .is_wysiwyg = "true";
defparam \regs[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \rfif.rdat2[2]~617 (
// Equation(s):
// \rfif.rdat2[2]~617_combout  = (\rfif.rdat2[2]~616_combout  & (((\regs[31][2]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[2]~616_combout  & (\regs[23][2]~q  & ((Instr_IF_18))))

	.dataa(\rfif.rdat2[2]~616_combout ),
	.datab(\regs[23][2]~q ),
	.datac(\regs[31][2]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~617_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~617 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[2]~617 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N21
dffeas \regs[29][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][2] .is_wysiwyg = "true";
defparam \regs[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N13
dffeas \regs[21][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][2] .is_wysiwyg = "true";
defparam \regs[21][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N31
dffeas \regs[17][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][2] .is_wysiwyg = "true";
defparam \regs[17][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N3
dffeas \regs[25][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][2] .is_wysiwyg = "true";
defparam \regs[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \rfif.rdat2[2]~609 (
// Equation(s):
// \rfif.rdat2[2]~609_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][2]~q ))) # (!Instr_IF_19 & (\regs[17][2]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[17][2]~q ),
	.datac(\regs[25][2]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~609_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~609 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[2]~609 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \rfif.rdat2[2]~610 (
// Equation(s):
// \rfif.rdat2[2]~610_combout  = (Instr_IF_18 & ((\rfif.rdat2[2]~609_combout  & (\regs[29][2]~q )) # (!\rfif.rdat2[2]~609_combout  & ((\regs[21][2]~q ))))) # (!Instr_IF_18 & (((\rfif.rdat2[2]~609_combout ))))

	.dataa(Instr_IF_18),
	.datab(\regs[29][2]~q ),
	.datac(\regs[21][2]~q ),
	.datad(\rfif.rdat2[2]~609_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~610_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~610 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[2]~610 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N31
dffeas \regs[16][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[16][2] .is_wysiwyg = "true";
defparam \regs[16][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N9
dffeas \regs[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][2] .is_wysiwyg = "true";
defparam \regs[20][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[2]~613 (
// Equation(s):
// \rfif.rdat2[2]~613_combout  = (Instr_IF_18 & ((Instr_IF_19) # ((\regs[20][2]~q )))) # (!Instr_IF_18 & (!Instr_IF_19 & (\regs[16][2]~q )))

	.dataa(Instr_IF_18),
	.datab(Instr_IF_19),
	.datac(\regs[16][2]~q ),
	.datad(\regs[20][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~613_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~613 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[2]~613 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N11
dffeas \regs[28][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][2] .is_wysiwyg = "true";
defparam \regs[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N29
dffeas \regs[24][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][2] .is_wysiwyg = "true";
defparam \regs[24][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \rfif.rdat2[2]~614 (
// Equation(s):
// \rfif.rdat2[2]~614_combout  = (Instr_IF_19 & ((\rfif.rdat2[2]~613_combout  & (\regs[28][2]~q )) # (!\rfif.rdat2[2]~613_combout  & ((\regs[24][2]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[2]~613_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[2]~613_combout ),
	.datac(\regs[28][2]~q ),
	.datad(\regs[24][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~614_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~614 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[2]~614 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N29
dffeas \regs[26][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][2] .is_wysiwyg = "true";
defparam \regs[26][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N7
dffeas \regs[30][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][2] .is_wysiwyg = "true";
defparam \regs[30][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N3
dffeas \regs[18][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][2] .is_wysiwyg = "true";
defparam \regs[18][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N13
dffeas \regs[22][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][2] .is_wysiwyg = "true";
defparam \regs[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[2]~611 (
// Equation(s):
// \rfif.rdat2[2]~611_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[22][2]~q ))) # (!Instr_IF_18 & (\regs[18][2]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[18][2]~q ),
	.datad(\regs[22][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~611_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~611 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[2]~611 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \rfif.rdat2[2]~612 (
// Equation(s):
// \rfif.rdat2[2]~612_combout  = (Instr_IF_19 & ((\rfif.rdat2[2]~611_combout  & ((\regs[30][2]~q ))) # (!\rfif.rdat2[2]~611_combout  & (\regs[26][2]~q )))) # (!Instr_IF_19 & (((\rfif.rdat2[2]~611_combout ))))

	.dataa(Instr_IF_19),
	.datab(\regs[26][2]~q ),
	.datac(\regs[30][2]~q ),
	.datad(\rfif.rdat2[2]~611_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~612_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~612 .lut_mask = 16'hF588;
defparam \rfif.rdat2[2]~612 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N10
cycloneive_lcell_comb \rfif.rdat2[2]~615 (
// Equation(s):
// \rfif.rdat2[2]~615_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & ((\rfif.rdat2[2]~612_combout ))) # (!Instr_IF_17 & (\rfif.rdat2[2]~614_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[2]~614_combout ),
	.datac(Instr_IF_17),
	.datad(\rfif.rdat2[2]~612_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~615_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~615 .lut_mask = 16'hF4A4;
defparam \rfif.rdat2[2]~615 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N0
cycloneive_lcell_comb \rfif.rdat2[2]~618 (
// Equation(s):
// \rfif.rdat2[2]~618_combout  = (Instr_IF_16 & ((\rfif.rdat2[2]~615_combout  & (\rfif.rdat2[2]~617_combout )) # (!\rfif.rdat2[2]~615_combout  & ((\rfif.rdat2[2]~610_combout ))))) # (!Instr_IF_16 & (((\rfif.rdat2[2]~615_combout ))))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[2]~617_combout ),
	.datac(\rfif.rdat2[2]~610_combout ),
	.datad(\rfif.rdat2[2]~615_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[2]~618_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[2]~618 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[2]~618 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \rfif.rdat1[2]~582 (
// Equation(s):
// \rfif.rdat1[2]~582_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][2]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[17][2]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[17][2]~q ),
	.datad(\regs[21][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~582_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~582 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[2]~582 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \rfif.rdat1[2]~583 (
// Equation(s):
// \rfif.rdat1[2]~583_combout  = (Instr_IF_24 & ((\rfif.rdat1[2]~582_combout  & ((\regs[29][2]~q ))) # (!\rfif.rdat1[2]~582_combout  & (\regs[25][2]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[2]~582_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[25][2]~q ),
	.datac(\regs[29][2]~q ),
	.datad(\rfif.rdat1[2]~582_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~583_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~583 .lut_mask = 16'hF588;
defparam \rfif.rdat1[2]~583 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N28
cycloneive_lcell_comb \rfif.rdat1[2]~584 (
// Equation(s):
// \rfif.rdat1[2]~584_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[24][2]~q ))) # (!Instr_IF_24 & (\regs[16][2]~q ))))

	.dataa(Instr_IF_23),
	.datab(\regs[16][2]~q ),
	.datac(\regs[24][2]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~584_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~584 .lut_mask = 16'hFA44;
defparam \rfif.rdat1[2]~584 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[2]~585 (
// Equation(s):
// \rfif.rdat1[2]~585_combout  = (Instr_IF_23 & ((\rfif.rdat1[2]~584_combout  & ((\regs[28][2]~q ))) # (!\rfif.rdat1[2]~584_combout  & (\regs[20][2]~q )))) # (!Instr_IF_23 & (\rfif.rdat1[2]~584_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[2]~584_combout ),
	.datac(\regs[20][2]~q ),
	.datad(\regs[28][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~585_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~585 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[2]~585 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \rfif.rdat1[2]~586 (
// Equation(s):
// \rfif.rdat1[2]~586_combout  = (Instr_IF_22 & (((Instr_IF_21)))) # (!Instr_IF_22 & ((Instr_IF_21 & (\rfif.rdat1[2]~583_combout )) # (!Instr_IF_21 & ((\rfif.rdat1[2]~585_combout )))))

	.dataa(Instr_IF_22),
	.datab(\rfif.rdat1[2]~583_combout ),
	.datac(Instr_IF_21),
	.datad(\rfif.rdat1[2]~585_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~586_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~586 .lut_mask = 16'hE5E0;
defparam \rfif.rdat1[2]~586 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[2]~587 (
// Equation(s):
// \rfif.rdat1[2]~587_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][2]~q ))) # (!Instr_IF_23 & (\regs[19][2]~q ))))

	.dataa(\regs[19][2]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[23][2]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~587_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~587 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[2]~587 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \regs[27][2]~feeder (
// Equation(s):
// \regs[27][2]~feeder_combout  = \input_a~129_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a12),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[27][2]~feeder .lut_mask = 16'hF0F0;
defparam \regs[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N11
dffeas \regs[27][2] (
	.clk(!CLK),
	.d(\regs[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][2] .is_wysiwyg = "true";
defparam \regs[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \rfif.rdat1[2]~588 (
// Equation(s):
// \rfif.rdat1[2]~588_combout  = (Instr_IF_24 & ((\rfif.rdat1[2]~587_combout  & (\regs[31][2]~q )) # (!\rfif.rdat1[2]~587_combout  & ((\regs[27][2]~q ))))) # (!Instr_IF_24 & (((\rfif.rdat1[2]~587_combout ))))

	.dataa(\regs[31][2]~q ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[2]~587_combout ),
	.datad(\regs[27][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~588_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~588 .lut_mask = 16'hBCB0;
defparam \rfif.rdat1[2]~588 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[2]~580 (
// Equation(s):
// \rfif.rdat1[2]~580_combout  = (Instr_IF_24 & (((\regs[26][2]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[18][2]~q  & ((!Instr_IF_23))))

	.dataa(\regs[18][2]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[26][2]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~580_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~580 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[2]~580 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[2]~581 (
// Equation(s):
// \rfif.rdat1[2]~581_combout  = (Instr_IF_23 & ((\rfif.rdat1[2]~580_combout  & (\regs[30][2]~q )) # (!\rfif.rdat1[2]~580_combout  & ((\regs[22][2]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[2]~580_combout ))))

	.dataa(Instr_IF_23),
	.datab(\regs[30][2]~q ),
	.datac(\regs[22][2]~q ),
	.datad(\rfif.rdat1[2]~580_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~581_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~581 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[2]~581 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \rfif.rdat1[2]~597 (
// Equation(s):
// \rfif.rdat1[2]~597_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][2]~q )) # (!Instr_IF_22 & ((\regs[12][2]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[14][2]~q ),
	.datad(\regs[12][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~597_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~597 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[2]~597 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N6
cycloneive_lcell_comb \rfif.rdat1[2]~598 (
// Equation(s):
// \rfif.rdat1[2]~598_combout  = (Instr_IF_21 & ((\rfif.rdat1[2]~597_combout  & (\regs[15][2]~q )) # (!\rfif.rdat1[2]~597_combout  & ((\regs[13][2]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[2]~597_combout ))))

	.dataa(\regs[15][2]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][2]~q ),
	.datad(\rfif.rdat1[2]~597_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~598_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~598 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[2]~598 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[2]~590 (
// Equation(s):
// \rfif.rdat1[2]~590_combout  = (Instr_IF_21 & (((\regs[9][2]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[8][2]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[8][2]~q ),
	.datac(\regs[9][2]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~590_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~590 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[2]~590 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \rfif.rdat1[2]~591 (
// Equation(s):
// \rfif.rdat1[2]~591_combout  = (Instr_IF_22 & ((\rfif.rdat1[2]~590_combout  & (\regs[11][2]~q )) # (!\rfif.rdat1[2]~590_combout  & ((\regs[10][2]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[2]~590_combout ))))

	.dataa(\regs[11][2]~q ),
	.datab(Instr_IF_22),
	.datac(\regs[10][2]~q ),
	.datad(\rfif.rdat1[2]~590_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~591_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~591 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[2]~591 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[2]~594 (
// Equation(s):
// \rfif.rdat1[2]~594_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & ((\regs[1][2]~q ))) # (!Instr_IF_21 & (\regs[0][2]~q ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[0][2]~q ),
	.datad(\regs[1][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~594_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~594 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[2]~594 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \rfif.rdat1[2]~595 (
// Equation(s):
// \rfif.rdat1[2]~595_combout  = (Instr_IF_22 & ((\rfif.rdat1[2]~594_combout  & ((\regs[3][2]~q ))) # (!\rfif.rdat1[2]~594_combout  & (\regs[2][2]~q )))) # (!Instr_IF_22 & (((\rfif.rdat1[2]~594_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[2][2]~q ),
	.datac(\rfif.rdat1[2]~594_combout ),
	.datad(\regs[3][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~595_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~595 .lut_mask = 16'hF858;
defparam \rfif.rdat1[2]~595 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N2
cycloneive_lcell_comb \rfif.rdat1[2]~592 (
// Equation(s):
// \rfif.rdat1[2]~592_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[6][2]~q ))) # (!Instr_IF_22 & (\regs[4][2]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[4][2]~q ),
	.datad(\regs[6][2]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~592_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~592 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[2]~592 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N21
dffeas \regs[7][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][2] .is_wysiwyg = "true";
defparam \regs[7][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \rfif.rdat1[2]~593 (
// Equation(s):
// \rfif.rdat1[2]~593_combout  = (\rfif.rdat1[2]~592_combout  & (((\regs[7][2]~q ) # (!Instr_IF_21)))) # (!\rfif.rdat1[2]~592_combout  & (\regs[5][2]~q  & ((Instr_IF_21))))

	.dataa(\regs[5][2]~q ),
	.datab(\rfif.rdat1[2]~592_combout ),
	.datac(\regs[7][2]~q ),
	.datad(Instr_IF_21),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~593_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~593 .lut_mask = 16'hE2CC;
defparam \rfif.rdat1[2]~593 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \rfif.rdat1[2]~596 (
// Equation(s):
// \rfif.rdat1[2]~596_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\rfif.rdat1[2]~593_combout )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\rfif.rdat1[2]~595_combout )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[2]~595_combout ),
	.datad(\rfif.rdat1[2]~593_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[2]~596_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[2]~596 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[2]~596 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N5
dffeas \regs[27][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][1] .is_wysiwyg = "true";
defparam \regs[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N27
dffeas \regs[31][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][1] .is_wysiwyg = "true";
defparam \regs[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \rfif.rdat2[1]~638 (
// Equation(s):
// \rfif.rdat2[1]~638_combout  = (\rfif.rdat2[1]~637_combout  & (((\regs[31][1]~q ) # (!Instr_IF_19)))) # (!\rfif.rdat2[1]~637_combout  & (\regs[27][1]~q  & ((Instr_IF_19))))

	.dataa(\rfif.rdat2[1]~637_combout ),
	.datab(\regs[27][1]~q ),
	.datac(\regs[31][1]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~638_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~638 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[1]~638 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N13
dffeas \regs[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][1] .is_wysiwyg = "true";
defparam \regs[22][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \regs[30][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][1] .is_wysiwyg = "true";
defparam \regs[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \rfif.rdat2[1]~631 (
// Equation(s):
// \rfif.rdat2[1]~631_combout  = (\rfif.rdat2[1]~630_combout  & (((\regs[30][1]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[1]~630_combout  & (Instr_IF_18 & (\regs[22][1]~q )))

	.dataa(\rfif.rdat2[1]~630_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[22][1]~q ),
	.datad(\regs[30][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~631_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~631 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[1]~631 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N3
dffeas \regs[28][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][1] .is_wysiwyg = "true";
defparam \regs[28][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N21
dffeas \regs[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][1] .is_wysiwyg = "true";
defparam \regs[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N2
cycloneive_lcell_comb \rfif.rdat2[1]~635 (
// Equation(s):
// \rfif.rdat2[1]~635_combout  = (\rfif.rdat2[1]~634_combout  & (((\regs[28][1]~q )) # (!Instr_IF_18))) # (!\rfif.rdat2[1]~634_combout  & (Instr_IF_18 & ((\regs[20][1]~q ))))

	.dataa(\rfif.rdat2[1]~634_combout ),
	.datab(Instr_IF_18),
	.datac(\regs[28][1]~q ),
	.datad(\regs[20][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~635_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~635 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[1]~635 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N11
dffeas \regs[17][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][1] .is_wysiwyg = "true";
defparam \regs[17][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N29
dffeas \regs[21][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][1] .is_wysiwyg = "true";
defparam \regs[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N10
cycloneive_lcell_comb \rfif.rdat2[1]~632 (
// Equation(s):
// \rfif.rdat2[1]~632_combout  = (Instr_IF_19 & (Instr_IF_18)) # (!Instr_IF_19 & ((Instr_IF_18 & ((\regs[21][1]~q ))) # (!Instr_IF_18 & (\regs[17][1]~q ))))

	.dataa(Instr_IF_19),
	.datab(Instr_IF_18),
	.datac(\regs[17][1]~q ),
	.datad(\regs[21][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~632_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~632 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[1]~632 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \regs[29][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][1] .is_wysiwyg = "true";
defparam \regs[29][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N29
dffeas \regs[25][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][1] .is_wysiwyg = "true";
defparam \regs[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \rfif.rdat2[1]~633 (
// Equation(s):
// \rfif.rdat2[1]~633_combout  = (Instr_IF_19 & ((\rfif.rdat2[1]~632_combout  & (\regs[29][1]~q )) # (!\rfif.rdat2[1]~632_combout  & ((\regs[25][1]~q ))))) # (!Instr_IF_19 & (\rfif.rdat2[1]~632_combout ))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[1]~632_combout ),
	.datac(\regs[29][1]~q ),
	.datad(\regs[25][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~633_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~633 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[1]~633 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[1]~636 (
// Equation(s):
// \rfif.rdat2[1]~636_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\rfif.rdat2[1]~633_combout ))) # (!Instr_IF_16 & (\rfif.rdat2[1]~635_combout ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\rfif.rdat2[1]~635_combout ),
	.datad(\rfif.rdat2[1]~633_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~636_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~636 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[1]~636 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N6
cycloneive_lcell_comb \rfif.rdat2[1]~639 (
// Equation(s):
// \rfif.rdat2[1]~639_combout  = (Instr_IF_17 & ((\rfif.rdat2[1]~636_combout  & (\rfif.rdat2[1]~638_combout )) # (!\rfif.rdat2[1]~636_combout  & ((\rfif.rdat2[1]~631_combout ))))) # (!Instr_IF_17 & (((\rfif.rdat2[1]~636_combout ))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[1]~638_combout ),
	.datac(\rfif.rdat2[1]~631_combout ),
	.datad(\rfif.rdat2[1]~636_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~639_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~639 .lut_mask = 16'hDDA0;
defparam \rfif.rdat2[1]~639 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N9
dffeas \regs[13][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][1] .is_wysiwyg = "true";
defparam \regs[13][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N15
dffeas \regs[15][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][1] .is_wysiwyg = "true";
defparam \regs[15][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N15
dffeas \regs[14][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][1] .is_wysiwyg = "true";
defparam \regs[14][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N25
dffeas \regs[12][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][1] .is_wysiwyg = "true";
defparam \regs[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N24
cycloneive_lcell_comb \rfif.rdat2[1]~647 (
// Equation(s):
// \rfif.rdat2[1]~647_combout  = (Instr_IF_17 & ((\regs[14][1]~q ) # ((Instr_IF_16)))) # (!Instr_IF_17 & (((\regs[12][1]~q  & !Instr_IF_16))))

	.dataa(Instr_IF_17),
	.datab(\regs[14][1]~q ),
	.datac(\regs[12][1]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~647_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~647 .lut_mask = 16'hAAD8;
defparam \rfif.rdat2[1]~647 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[1]~648 (
// Equation(s):
// \rfif.rdat2[1]~648_combout  = (Instr_IF_16 & ((\rfif.rdat2[1]~647_combout  & ((\regs[15][1]~q ))) # (!\rfif.rdat2[1]~647_combout  & (\regs[13][1]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[1]~647_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[13][1]~q ),
	.datac(\regs[15][1]~q ),
	.datad(\rfif.rdat2[1]~647_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~648_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~648 .lut_mask = 16'hF588;
defparam \rfif.rdat2[1]~648 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N9
dffeas \regs[5][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][1] .is_wysiwyg = "true";
defparam \regs[5][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N23
dffeas \regs[7][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][1] .is_wysiwyg = "true";
defparam \regs[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N5
dffeas \regs[6][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][1] .is_wysiwyg = "true";
defparam \regs[6][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N15
dffeas \regs[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][1] .is_wysiwyg = "true";
defparam \regs[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \rfif.rdat2[1]~642 (
// Equation(s):
// \rfif.rdat2[1]~642_combout  = (Instr_IF_16 & (((Instr_IF_17)))) # (!Instr_IF_16 & ((Instr_IF_17 & (\regs[6][1]~q )) # (!Instr_IF_17 & ((\regs[4][1]~q )))))

	.dataa(Instr_IF_16),
	.datab(\regs[6][1]~q ),
	.datac(\regs[4][1]~q ),
	.datad(Instr_IF_17),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~642_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~642 .lut_mask = 16'hEE50;
defparam \rfif.rdat2[1]~642 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \rfif.rdat2[1]~643 (
// Equation(s):
// \rfif.rdat2[1]~643_combout  = (Instr_IF_16 & ((\rfif.rdat2[1]~642_combout  & ((\regs[7][1]~q ))) # (!\rfif.rdat2[1]~642_combout  & (\regs[5][1]~q )))) # (!Instr_IF_16 & (((\rfif.rdat2[1]~642_combout ))))

	.dataa(Instr_IF_16),
	.datab(\regs[5][1]~q ),
	.datac(\regs[7][1]~q ),
	.datad(\rfif.rdat2[1]~642_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~643_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~643 .lut_mask = 16'hF588;
defparam \rfif.rdat2[1]~643 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \regs[2][1]~feeder (
// Equation(s):
// \regs[2][1]~feeder_combout  = \input_a~132_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(input_a13),
	.datad(gnd),
	.cin(gnd),
	.combout(\regs[2][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[2][1]~feeder .lut_mask = 16'hF0F0;
defparam \regs[2][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N5
dffeas \regs[2][1] (
	.clk(!CLK),
	.d(\regs[2][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][1] .is_wysiwyg = "true";
defparam \regs[2][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N15
dffeas \regs[3][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][1] .is_wysiwyg = "true";
defparam \regs[3][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N31
dffeas \regs[0][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][1] .is_wysiwyg = "true";
defparam \regs[0][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N9
dffeas \regs[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][1] .is_wysiwyg = "true";
defparam \regs[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[1]~644 (
// Equation(s):
// \rfif.rdat2[1]~644_combout  = (Instr_IF_16 & ((Instr_IF_17) # ((\regs[1][1]~q )))) # (!Instr_IF_16 & (!Instr_IF_17 & (\regs[0][1]~q )))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][1]~q ),
	.datad(\regs[1][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~644_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~644 .lut_mask = 16'hBA98;
defparam \rfif.rdat2[1]~644 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \rfif.rdat2[1]~645 (
// Equation(s):
// \rfif.rdat2[1]~645_combout  = (Instr_IF_17 & ((\rfif.rdat2[1]~644_combout  & ((\regs[3][1]~q ))) # (!\rfif.rdat2[1]~644_combout  & (\regs[2][1]~q )))) # (!Instr_IF_17 & (((\rfif.rdat2[1]~644_combout ))))

	.dataa(Instr_IF_17),
	.datab(\regs[2][1]~q ),
	.datac(\regs[3][1]~q ),
	.datad(\rfif.rdat2[1]~644_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~645_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~645 .lut_mask = 16'hF588;
defparam \rfif.rdat2[1]~645 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N30
cycloneive_lcell_comb \rfif.rdat2[1]~646 (
// Equation(s):
// \rfif.rdat2[1]~646_combout  = (Instr_IF_18 & ((\rfif.rdat2[1]~643_combout ) # ((Instr_IF_19)))) # (!Instr_IF_18 & (((!Instr_IF_19 & \rfif.rdat2[1]~645_combout ))))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[1]~643_combout ),
	.datac(Instr_IF_19),
	.datad(\rfif.rdat2[1]~645_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~646_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~646 .lut_mask = 16'hADA8;
defparam \rfif.rdat2[1]~646 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N21
dffeas \regs[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][1] .is_wysiwyg = "true";
defparam \regs[10][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N5
dffeas \regs[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][1] .is_wysiwyg = "true";
defparam \regs[9][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N4
cycloneive_lcell_comb \rfif.rdat2[1]~640 (
// Equation(s):
// \rfif.rdat2[1]~640_combout  = (Instr_IF_17 & (((Instr_IF_16)))) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[9][1]~q ))) # (!Instr_IF_16 & (\regs[8][1]~q ))))

	.dataa(\regs[8][1]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[9][1]~q ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~640_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~640 .lut_mask = 16'hFC22;
defparam \rfif.rdat2[1]~640 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N20
cycloneive_lcell_comb \rfif.rdat2[1]~641 (
// Equation(s):
// \rfif.rdat2[1]~641_combout  = (Instr_IF_17 & ((\rfif.rdat2[1]~640_combout  & (\regs[11][1]~q )) # (!\rfif.rdat2[1]~640_combout  & ((\regs[10][1]~q ))))) # (!Instr_IF_17 & (((\rfif.rdat2[1]~640_combout ))))

	.dataa(\regs[11][1]~q ),
	.datab(Instr_IF_17),
	.datac(\regs[10][1]~q ),
	.datad(\rfif.rdat2[1]~640_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~641_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~641 .lut_mask = 16'hBBC0;
defparam \rfif.rdat2[1]~641 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N8
cycloneive_lcell_comb \rfif.rdat2[1]~649 (
// Equation(s):
// \rfif.rdat2[1]~649_combout  = (Instr_IF_19 & ((\rfif.rdat2[1]~646_combout  & (\rfif.rdat2[1]~648_combout )) # (!\rfif.rdat2[1]~646_combout  & ((\rfif.rdat2[1]~641_combout ))))) # (!Instr_IF_19 & (((\rfif.rdat2[1]~646_combout ))))

	.dataa(Instr_IF_19),
	.datab(\rfif.rdat2[1]~648_combout ),
	.datac(\rfif.rdat2[1]~646_combout ),
	.datad(\rfif.rdat2[1]~641_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[1]~649_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[1]~649 .lut_mask = 16'hDAD0;
defparam \rfif.rdat2[1]~649 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \regs[26][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][1] .is_wysiwyg = "true";
defparam \regs[26][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N7
dffeas \regs[18][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][1] .is_wysiwyg = "true";
defparam \regs[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \rfif.rdat1[1]~602 (
// Equation(s):
// \rfif.rdat1[1]~602_combout  = (Instr_IF_24 & (Instr_IF_23)) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[22][1]~q ))) # (!Instr_IF_23 & (\regs[18][1]~q ))))

	.dataa(Instr_IF_24),
	.datab(Instr_IF_23),
	.datac(\regs[18][1]~q ),
	.datad(\regs[22][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~602_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~602 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[1]~602 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \rfif.rdat1[1]~603 (
// Equation(s):
// \rfif.rdat1[1]~603_combout  = (Instr_IF_24 & ((\rfif.rdat1[1]~602_combout  & ((\regs[30][1]~q ))) # (!\rfif.rdat1[1]~602_combout  & (\regs[26][1]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[1]~602_combout ))))

	.dataa(Instr_IF_24),
	.datab(\regs[26][1]~q ),
	.datac(\regs[30][1]~q ),
	.datad(\rfif.rdat1[1]~602_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~603_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~603 .lut_mask = 16'hF588;
defparam \rfif.rdat1[1]~603 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N20
cycloneive_lcell_comb \rfif.rdat1[1]~604 (
// Equation(s):
// \rfif.rdat1[1]~604_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[20][1]~q ))) # (!Instr_IF_23 & (\regs[16][1]~q ))))

	.dataa(\regs[16][1]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[20][1]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~604_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~604 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[1]~604 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N13
dffeas \regs[24][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][1] .is_wysiwyg = "true";
defparam \regs[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[1]~605 (
// Equation(s):
// \rfif.rdat1[1]~605_combout  = (\rfif.rdat1[1]~604_combout  & ((\regs[28][1]~q ) # ((!Instr_IF_24)))) # (!\rfif.rdat1[1]~604_combout  & (((\regs[24][1]~q  & Instr_IF_24))))

	.dataa(\regs[28][1]~q ),
	.datab(\rfif.rdat1[1]~604_combout ),
	.datac(\regs[24][1]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~605_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~605 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[1]~605 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \rfif.rdat1[1]~606 (
// Equation(s):
// \rfif.rdat1[1]~606_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\rfif.rdat1[1]~603_combout )))) # (!Instr_IF_22 & (!Instr_IF_21 & ((\rfif.rdat1[1]~605_combout ))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\rfif.rdat1[1]~603_combout ),
	.datad(\rfif.rdat1[1]~605_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~606_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~606 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[1]~606 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N15
dffeas \regs[19][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[19][1] .is_wysiwyg = "true";
defparam \regs[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \rfif.rdat1[1]~607 (
// Equation(s):
// \rfif.rdat1[1]~607_combout  = (Instr_IF_24 & (((\regs[27][1]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[19][1]~q  & ((!Instr_IF_23))))

	.dataa(Instr_IF_24),
	.datab(\regs[19][1]~q ),
	.datac(\regs[27][1]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~607_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~607 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[1]~607 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N21
dffeas \regs[23][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][1] .is_wysiwyg = "true";
defparam \regs[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[1]~608 (
// Equation(s):
// \rfif.rdat1[1]~608_combout  = (Instr_IF_23 & ((\rfif.rdat1[1]~607_combout  & ((\regs[31][1]~q ))) # (!\rfif.rdat1[1]~607_combout  & (\regs[23][1]~q )))) # (!Instr_IF_23 & (\rfif.rdat1[1]~607_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[1]~607_combout ),
	.datac(\regs[23][1]~q ),
	.datad(\regs[31][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~608_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~608 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[1]~608 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \rfif.rdat1[1]~600 (
// Equation(s):
// \rfif.rdat1[1]~600_combout  = (Instr_IF_23 & (((Instr_IF_24)))) # (!Instr_IF_23 & ((Instr_IF_24 & ((\regs[25][1]~q ))) # (!Instr_IF_24 & (\regs[17][1]~q ))))

	.dataa(\regs[17][1]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[25][1]~q ),
	.datad(Instr_IF_24),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~600_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~600 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[1]~600 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N28
cycloneive_lcell_comb \rfif.rdat1[1]~601 (
// Equation(s):
// \rfif.rdat1[1]~601_combout  = (Instr_IF_23 & ((\rfif.rdat1[1]~600_combout  & (\regs[29][1]~q )) # (!\rfif.rdat1[1]~600_combout  & ((\regs[21][1]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[1]~600_combout ))))

	.dataa(\regs[29][1]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[21][1]~q ),
	.datad(\rfif.rdat1[1]~600_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~601_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~601 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[1]~601 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \rfif.rdat1[1]~614 (
// Equation(s):
// \rfif.rdat1[1]~614_combout  = (Instr_IF_21 & (((Instr_IF_22)))) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[2][1]~q ))) # (!Instr_IF_22 & (\regs[0][1]~q ))))

	.dataa(\regs[0][1]~q ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\regs[2][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~614_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~614 .lut_mask = 16'hF2C2;
defparam \rfif.rdat1[1]~614 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \rfif.rdat1[1]~615 (
// Equation(s):
// \rfif.rdat1[1]~615_combout  = (Instr_IF_21 & ((\rfif.rdat1[1]~614_combout  & (\regs[3][1]~q )) # (!\rfif.rdat1[1]~614_combout  & ((\regs[1][1]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[1]~614_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[3][1]~q ),
	.datac(\regs[1][1]~q ),
	.datad(\rfif.rdat1[1]~614_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~615_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~615 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[1]~615 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N3
dffeas \regs[11][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][1] .is_wysiwyg = "true";
defparam \regs[11][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N15
dffeas \regs[8][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][1] .is_wysiwyg = "true";
defparam \regs[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N14
cycloneive_lcell_comb \rfif.rdat1[1]~612 (
// Equation(s):
// \rfif.rdat1[1]~612_combout  = (Instr_IF_22 & ((Instr_IF_21) # ((\regs[10][1]~q )))) # (!Instr_IF_22 & (!Instr_IF_21 & (\regs[8][1]~q )))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[8][1]~q ),
	.datad(\regs[10][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~612_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~612 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[1]~612 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N2
cycloneive_lcell_comb \rfif.rdat1[1]~613 (
// Equation(s):
// \rfif.rdat1[1]~613_combout  = (Instr_IF_21 & ((\rfif.rdat1[1]~612_combout  & ((\regs[11][1]~q ))) # (!\rfif.rdat1[1]~612_combout  & (\regs[9][1]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[1]~612_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[9][1]~q ),
	.datac(\regs[11][1]~q ),
	.datad(\rfif.rdat1[1]~612_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~613_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~613 .lut_mask = 16'hF588;
defparam \rfif.rdat1[1]~613 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[1]~616 (
// Equation(s):
// \rfif.rdat1[1]~616_combout  = (Instr_IF_24 & (((\rfif.rdat1[1]~613_combout ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\rfif.rdat1[1]~615_combout  & ((!Instr_IF_23))))

	.dataa(\rfif.rdat1[1]~615_combout ),
	.datab(\rfif.rdat1[1]~613_combout ),
	.datac(Instr_IF_24),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~616_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~616 .lut_mask = 16'hF0CA;
defparam \rfif.rdat1[1]~616 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[1]~617 (
// Equation(s):
// \rfif.rdat1[1]~617_combout  = (Instr_IF_21 & ((Instr_IF_22) # ((\regs[13][1]~q )))) # (!Instr_IF_21 & (!Instr_IF_22 & ((\regs[12][1]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[13][1]~q ),
	.datad(\regs[12][1]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~617_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~617 .lut_mask = 16'hB9A8;
defparam \rfif.rdat1[1]~617 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \rfif.rdat1[1]~618 (
// Equation(s):
// \rfif.rdat1[1]~618_combout  = (\rfif.rdat1[1]~617_combout  & ((\regs[15][1]~q ) # ((!Instr_IF_22)))) # (!\rfif.rdat1[1]~617_combout  & (((\regs[14][1]~q  & Instr_IF_22))))

	.dataa(\regs[15][1]~q ),
	.datab(\rfif.rdat1[1]~617_combout ),
	.datac(\regs[14][1]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~618_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~618 .lut_mask = 16'hB8CC;
defparam \rfif.rdat1[1]~618 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \rfif.rdat1[1]~610 (
// Equation(s):
// \rfif.rdat1[1]~610_combout  = (Instr_IF_21 & (((\regs[5][1]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[4][1]~q  & ((!Instr_IF_22))))

	.dataa(\regs[4][1]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[5][1]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~610_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~610 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[1]~610 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \rfif.rdat1[1]~611 (
// Equation(s):
// \rfif.rdat1[1]~611_combout  = (Instr_IF_22 & ((\rfif.rdat1[1]~610_combout  & (\regs[7][1]~q )) # (!\rfif.rdat1[1]~610_combout  & ((\regs[6][1]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[1]~610_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[7][1]~q ),
	.datac(\regs[6][1]~q ),
	.datad(\rfif.rdat1[1]~610_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[1]~611_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[1]~611 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[1]~611 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N9
dffeas \regs[0][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[0][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[0][0] .is_wysiwyg = "true";
defparam \regs[0][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N19
dffeas \regs[2][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[2][0] .is_wysiwyg = "true";
defparam \regs[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \rfif.rdat2[0]~665 (
// Equation(s):
// \rfif.rdat2[0]~665_combout  = (Instr_IF_16 & (Instr_IF_17)) # (!Instr_IF_16 & ((Instr_IF_17 & ((\regs[2][0]~q ))) # (!Instr_IF_17 & (\regs[0][0]~q ))))

	.dataa(Instr_IF_16),
	.datab(Instr_IF_17),
	.datac(\regs[0][0]~q ),
	.datad(\regs[2][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~665_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~665 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[0]~665 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N31
dffeas \regs[3][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[3][0] .is_wysiwyg = "true";
defparam \regs[3][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N25
dffeas \regs[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[1][0] .is_wysiwyg = "true";
defparam \regs[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \rfif.rdat2[0]~666 (
// Equation(s):
// \rfif.rdat2[0]~666_combout  = (Instr_IF_16 & ((\rfif.rdat2[0]~665_combout  & (\regs[3][0]~q )) # (!\rfif.rdat2[0]~665_combout  & ((\regs[1][0]~q ))))) # (!Instr_IF_16 & (\rfif.rdat2[0]~665_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[0]~665_combout ),
	.datac(\regs[3][0]~q ),
	.datad(\regs[1][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~666_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~666 .lut_mask = 16'hE6C4;
defparam \rfif.rdat2[0]~666 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \rfif.rdat2[0]~667 (
// Equation(s):
// \rfif.rdat2[0]~667_combout  = (Instr_IF_19 & ((\rfif.rdat2[0]~664_combout ) # ((Instr_IF_18)))) # (!Instr_IF_19 & (((\rfif.rdat2[0]~666_combout  & !Instr_IF_18))))

	.dataa(\rfif.rdat2[0]~664_combout ),
	.datab(Instr_IF_19),
	.datac(\rfif.rdat2[0]~666_combout ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~667_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~667 .lut_mask = 16'hCCB8;
defparam \rfif.rdat2[0]~667 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N27
dffeas \regs[12][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[12][0] .is_wysiwyg = "true";
defparam \regs[12][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N23
dffeas \regs[13][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[13][0] .is_wysiwyg = "true";
defparam \regs[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \rfif.rdat2[0]~668 (
// Equation(s):
// \rfif.rdat2[0]~668_combout  = (Instr_IF_17 & (Instr_IF_16)) # (!Instr_IF_17 & ((Instr_IF_16 & ((\regs[13][0]~q ))) # (!Instr_IF_16 & (\regs[12][0]~q ))))

	.dataa(Instr_IF_17),
	.datab(Instr_IF_16),
	.datac(\regs[12][0]~q ),
	.datad(\regs[13][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~668_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~668 .lut_mask = 16'hDC98;
defparam \rfif.rdat2[0]~668 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \regs[15][0]~feeder (
// Equation(s):
// \regs[15][0]~feeder_combout  = \input_a~135_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(input_a14),
	.cin(gnd),
	.combout(\regs[15][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \regs[15][0]~feeder .lut_mask = 16'hFF00;
defparam \regs[15][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N3
dffeas \regs[15][0] (
	.clk(!CLK),
	.d(\regs[15][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[15][0] .is_wysiwyg = "true";
defparam \regs[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \rfif.rdat2[0]~669 (
// Equation(s):
// \rfif.rdat2[0]~669_combout  = (\rfif.rdat2[0]~668_combout  & (((\regs[15][0]~q ) # (!Instr_IF_17)))) # (!\rfif.rdat2[0]~668_combout  & (\regs[14][0]~q  & (Instr_IF_17)))

	.dataa(\regs[14][0]~q ),
	.datab(\rfif.rdat2[0]~668_combout ),
	.datac(Instr_IF_17),
	.datad(\regs[15][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~669_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~669 .lut_mask = 16'hEC2C;
defparam \rfif.rdat2[0]~669 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N13
dffeas \regs[6][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[6][0] .is_wysiwyg = "true";
defparam \regs[6][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N5
dffeas \regs[7][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[7][0] .is_wysiwyg = "true";
defparam \regs[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \rfif.rdat2[0]~662 (
// Equation(s):
// \rfif.rdat2[0]~662_combout  = (\rfif.rdat2[0]~661_combout  & (((\regs[7][0]~q )) # (!Instr_IF_17))) # (!\rfif.rdat2[0]~661_combout  & (Instr_IF_17 & (\regs[6][0]~q )))

	.dataa(\rfif.rdat2[0]~661_combout ),
	.datab(Instr_IF_17),
	.datac(\regs[6][0]~q ),
	.datad(\regs[7][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~662_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~662 .lut_mask = 16'hEA62;
defparam \rfif.rdat2[0]~662 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \rfif.rdat2[0]~670 (
// Equation(s):
// \rfif.rdat2[0]~670_combout  = (\rfif.rdat2[0]~667_combout  & ((\rfif.rdat2[0]~669_combout ) # ((!Instr_IF_18)))) # (!\rfif.rdat2[0]~667_combout  & (((\rfif.rdat2[0]~662_combout  & Instr_IF_18))))

	.dataa(\rfif.rdat2[0]~667_combout ),
	.datab(\rfif.rdat2[0]~669_combout ),
	.datac(\rfif.rdat2[0]~662_combout ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~670_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~670 .lut_mask = 16'hD8AA;
defparam \rfif.rdat2[0]~670 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N7
dffeas \regs[28][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[28][0] .is_wysiwyg = "true";
defparam \regs[28][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N9
dffeas \regs[24][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[24][0] .is_wysiwyg = "true";
defparam \regs[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N6
cycloneive_lcell_comb \rfif.rdat2[0]~656 (
// Equation(s):
// \rfif.rdat2[0]~656_combout  = (\rfif.rdat2[0]~655_combout  & (((\regs[28][0]~q )) # (!Instr_IF_19))) # (!\rfif.rdat2[0]~655_combout  & (Instr_IF_19 & ((\regs[24][0]~q ))))

	.dataa(\rfif.rdat2[0]~655_combout ),
	.datab(Instr_IF_19),
	.datac(\regs[28][0]~q ),
	.datad(\regs[24][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~656_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~656 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[0]~656 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N27
dffeas \regs[30][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[30][0] .is_wysiwyg = "true";
defparam \regs[30][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N1
dffeas \regs[26][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[26][0] .is_wysiwyg = "true";
defparam \regs[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \rfif.rdat2[0]~654 (
// Equation(s):
// \rfif.rdat2[0]~654_combout  = (\rfif.rdat2[0]~653_combout  & (((\regs[30][0]~q )) # (!Instr_IF_19))) # (!\rfif.rdat2[0]~653_combout  & (Instr_IF_19 & ((\regs[26][0]~q ))))

	.dataa(\rfif.rdat2[0]~653_combout ),
	.datab(Instr_IF_19),
	.datac(\regs[30][0]~q ),
	.datad(\regs[26][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~654_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~654 .lut_mask = 16'hE6A2;
defparam \rfif.rdat2[0]~654 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \rfif.rdat2[0]~657 (
// Equation(s):
// \rfif.rdat2[0]~657_combout  = (Instr_IF_17 & (((\rfif.rdat2[0]~654_combout ) # (Instr_IF_16)))) # (!Instr_IF_17 & (\rfif.rdat2[0]~656_combout  & ((!Instr_IF_16))))

	.dataa(Instr_IF_17),
	.datab(\rfif.rdat2[0]~656_combout ),
	.datac(\rfif.rdat2[0]~654_combout ),
	.datad(Instr_IF_16),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~657_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~657 .lut_mask = 16'hAAE4;
defparam \rfif.rdat2[0]~657 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N11
dffeas \regs[17][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[17][0] .is_wysiwyg = "true";
defparam \regs[17][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N23
dffeas \regs[25][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[25][0] .is_wysiwyg = "true";
defparam \regs[25][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \rfif.rdat2[0]~651 (
// Equation(s):
// \rfif.rdat2[0]~651_combout  = (Instr_IF_18 & (((Instr_IF_19)))) # (!Instr_IF_18 & ((Instr_IF_19 & ((\regs[25][0]~q ))) # (!Instr_IF_19 & (\regs[17][0]~q ))))

	.dataa(Instr_IF_18),
	.datab(\regs[17][0]~q ),
	.datac(\regs[25][0]~q ),
	.datad(Instr_IF_19),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~651_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~651 .lut_mask = 16'hFA44;
defparam \rfif.rdat2[0]~651 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N17
dffeas \regs[21][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[21][0] .is_wysiwyg = "true";
defparam \regs[21][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \regs[29][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[29][0] .is_wysiwyg = "true";
defparam \regs[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \rfif.rdat2[0]~652 (
// Equation(s):
// \rfif.rdat2[0]~652_combout  = (Instr_IF_18 & ((\rfif.rdat2[0]~651_combout  & ((\regs[29][0]~q ))) # (!\rfif.rdat2[0]~651_combout  & (\regs[21][0]~q )))) # (!Instr_IF_18 & (\rfif.rdat2[0]~651_combout ))

	.dataa(Instr_IF_18),
	.datab(\rfif.rdat2[0]~651_combout ),
	.datac(\regs[21][0]~q ),
	.datad(\regs[29][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~652_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~652 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[0]~652 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N1
dffeas \regs[23][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[23][0] .is_wysiwyg = "true";
defparam \regs[23][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \regs[31][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[31][0] .is_wysiwyg = "true";
defparam \regs[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \rfif.rdat2[0]~659 (
// Equation(s):
// \rfif.rdat2[0]~659_combout  = (\rfif.rdat2[0]~658_combout  & (((\regs[31][0]~q ) # (!Instr_IF_18)))) # (!\rfif.rdat2[0]~658_combout  & (\regs[23][0]~q  & ((Instr_IF_18))))

	.dataa(\rfif.rdat2[0]~658_combout ),
	.datab(\regs[23][0]~q ),
	.datac(\regs[31][0]~q ),
	.datad(Instr_IF_18),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~659_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~659 .lut_mask = 16'hE4AA;
defparam \rfif.rdat2[0]~659 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \rfif.rdat2[0]~660 (
// Equation(s):
// \rfif.rdat2[0]~660_combout  = (Instr_IF_16 & ((\rfif.rdat2[0]~657_combout  & ((\rfif.rdat2[0]~659_combout ))) # (!\rfif.rdat2[0]~657_combout  & (\rfif.rdat2[0]~652_combout )))) # (!Instr_IF_16 & (\rfif.rdat2[0]~657_combout ))

	.dataa(Instr_IF_16),
	.datab(\rfif.rdat2[0]~657_combout ),
	.datac(\rfif.rdat2[0]~652_combout ),
	.datad(\rfif.rdat2[0]~659_combout ),
	.cin(gnd),
	.combout(\rfif.rdat2[0]~660_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat2[0]~660 .lut_mask = 16'hEC64;
defparam \rfif.rdat2[0]~660 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N29
dffeas \regs[22][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[22][0] .is_wysiwyg = "true";
defparam \regs[22][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N11
dffeas \regs[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[18][0] .is_wysiwyg = "true";
defparam \regs[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \rfif.rdat1[0]~620 (
// Equation(s):
// \rfif.rdat1[0]~620_combout  = (Instr_IF_23 & (Instr_IF_24)) # (!Instr_IF_23 & ((Instr_IF_24 & (\regs[26][0]~q )) # (!Instr_IF_24 & ((\regs[18][0]~q )))))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[26][0]~q ),
	.datad(\regs[18][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~620_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~620 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[0]~620 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \rfif.rdat1[0]~621 (
// Equation(s):
// \rfif.rdat1[0]~621_combout  = (Instr_IF_23 & ((\rfif.rdat1[0]~620_combout  & (\regs[30][0]~q )) # (!\rfif.rdat1[0]~620_combout  & ((\regs[22][0]~q ))))) # (!Instr_IF_23 & (((\rfif.rdat1[0]~620_combout ))))

	.dataa(\regs[30][0]~q ),
	.datab(Instr_IF_23),
	.datac(\regs[22][0]~q ),
	.datad(\rfif.rdat1[0]~620_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~621_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~621 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[0]~621 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \rfif.rdat1[0]~627 (
// Equation(s):
// \rfif.rdat1[0]~627_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\regs[23][0]~q ))) # (!Instr_IF_23 & (\regs[19][0]~q ))))

	.dataa(\regs[19][0]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[23][0]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~627_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~627 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[0]~627 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N21
dffeas \regs[27][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[27][0] .is_wysiwyg = "true";
defparam \regs[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \rfif.rdat1[0]~628 (
// Equation(s):
// \rfif.rdat1[0]~628_combout  = (Instr_IF_24 & ((\rfif.rdat1[0]~627_combout  & ((\regs[31][0]~q ))) # (!\rfif.rdat1[0]~627_combout  & (\regs[27][0]~q )))) # (!Instr_IF_24 & (\rfif.rdat1[0]~627_combout ))

	.dataa(Instr_IF_24),
	.datab(\rfif.rdat1[0]~627_combout ),
	.datac(\regs[27][0]~q ),
	.datad(\regs[31][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~628_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~628 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[0]~628 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \rfif.rdat1[0]~622 (
// Equation(s):
// \rfif.rdat1[0]~622_combout  = (Instr_IF_23 & ((Instr_IF_24) # ((\regs[21][0]~q )))) # (!Instr_IF_23 & (!Instr_IF_24 & (\regs[17][0]~q )))

	.dataa(Instr_IF_23),
	.datab(Instr_IF_24),
	.datac(\regs[17][0]~q ),
	.datad(\regs[21][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~622_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~622 .lut_mask = 16'hBA98;
defparam \rfif.rdat1[0]~622 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[0]~623 (
// Equation(s):
// \rfif.rdat1[0]~623_combout  = (Instr_IF_24 & ((\rfif.rdat1[0]~622_combout  & ((\regs[29][0]~q ))) # (!\rfif.rdat1[0]~622_combout  & (\regs[25][0]~q )))) # (!Instr_IF_24 & (((\rfif.rdat1[0]~622_combout ))))

	.dataa(\regs[25][0]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[29][0]~q ),
	.datad(\rfif.rdat1[0]~622_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~623_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~623 .lut_mask = 16'hF388;
defparam \rfif.rdat1[0]~623 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N8
cycloneive_lcell_comb \rfif.rdat1[0]~624 (
// Equation(s):
// \rfif.rdat1[0]~624_combout  = (Instr_IF_24 & (((\regs[24][0]~q ) # (Instr_IF_23)))) # (!Instr_IF_24 & (\regs[16][0]~q  & ((!Instr_IF_23))))

	.dataa(\regs[16][0]~q ),
	.datab(Instr_IF_24),
	.datac(\regs[24][0]~q ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~624_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~624 .lut_mask = 16'hCCE2;
defparam \rfif.rdat1[0]~624 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N17
dffeas \regs[20][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[20][0] .is_wysiwyg = "true";
defparam \regs[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N16
cycloneive_lcell_comb \rfif.rdat1[0]~625 (
// Equation(s):
// \rfif.rdat1[0]~625_combout  = (Instr_IF_23 & ((\rfif.rdat1[0]~624_combout  & ((\regs[28][0]~q ))) # (!\rfif.rdat1[0]~624_combout  & (\regs[20][0]~q )))) # (!Instr_IF_23 & (\rfif.rdat1[0]~624_combout ))

	.dataa(Instr_IF_23),
	.datab(\rfif.rdat1[0]~624_combout ),
	.datac(\regs[20][0]~q ),
	.datad(\regs[28][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~625_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~625 .lut_mask = 16'hEC64;
defparam \rfif.rdat1[0]~625 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \rfif.rdat1[0]~626 (
// Equation(s):
// \rfif.rdat1[0]~626_combout  = (Instr_IF_21 & ((\rfif.rdat1[0]~623_combout ) # ((Instr_IF_22)))) # (!Instr_IF_21 & (((!Instr_IF_22 & \rfif.rdat1[0]~625_combout ))))

	.dataa(\rfif.rdat1[0]~623_combout ),
	.datab(Instr_IF_21),
	.datac(Instr_IF_22),
	.datad(\rfif.rdat1[0]~625_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~626_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~626 .lut_mask = 16'hCBC8;
defparam \rfif.rdat1[0]~626 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N23
dffeas \regs[8][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[8][0] .is_wysiwyg = "true";
defparam \regs[8][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N17
dffeas \regs[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[9][0] .is_wysiwyg = "true";
defparam \regs[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \rfif.rdat1[0]~630 (
// Equation(s):
// \rfif.rdat1[0]~630_combout  = (Instr_IF_21 & (((\regs[9][0]~q ) # (Instr_IF_22)))) # (!Instr_IF_21 & (\regs[8][0]~q  & ((!Instr_IF_22))))

	.dataa(Instr_IF_21),
	.datab(\regs[8][0]~q ),
	.datac(\regs[9][0]~q ),
	.datad(Instr_IF_22),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~630_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~630 .lut_mask = 16'hAAE4;
defparam \rfif.rdat1[0]~630 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N29
dffeas \regs[10][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[10][0] .is_wysiwyg = "true";
defparam \regs[10][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N23
dffeas \regs[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[11][0] .is_wysiwyg = "true";
defparam \regs[11][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \rfif.rdat1[0]~631 (
// Equation(s):
// \rfif.rdat1[0]~631_combout  = (\rfif.rdat1[0]~630_combout  & (((\regs[11][0]~q )) # (!Instr_IF_22))) # (!\rfif.rdat1[0]~630_combout  & (Instr_IF_22 & (\regs[10][0]~q )))

	.dataa(\rfif.rdat1[0]~630_combout ),
	.datab(Instr_IF_22),
	.datac(\regs[10][0]~q ),
	.datad(\regs[11][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~631_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~631 .lut_mask = 16'hEA62;
defparam \rfif.rdat1[0]~631 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N25
dffeas \regs[14][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[14][0] .is_wysiwyg = "true";
defparam \regs[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N24
cycloneive_lcell_comb \rfif.rdat1[0]~637 (
// Equation(s):
// \rfif.rdat1[0]~637_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & (\regs[14][0]~q )) # (!Instr_IF_22 & ((\regs[12][0]~q )))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[14][0]~q ),
	.datad(\regs[12][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~637_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~637 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[0]~637 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \rfif.rdat1[0]~638 (
// Equation(s):
// \rfif.rdat1[0]~638_combout  = (Instr_IF_21 & ((\rfif.rdat1[0]~637_combout  & (\regs[15][0]~q )) # (!\rfif.rdat1[0]~637_combout  & ((\regs[13][0]~q ))))) # (!Instr_IF_21 & (((\rfif.rdat1[0]~637_combout ))))

	.dataa(\regs[15][0]~q ),
	.datab(Instr_IF_21),
	.datac(\regs[13][0]~q ),
	.datad(\rfif.rdat1[0]~637_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~638_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~638 .lut_mask = 16'hBBC0;
defparam \rfif.rdat1[0]~638 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \rfif.rdat1[0]~634 (
// Equation(s):
// \rfif.rdat1[0]~634_combout  = (Instr_IF_22 & (Instr_IF_21)) # (!Instr_IF_22 & ((Instr_IF_21 & (\regs[1][0]~q )) # (!Instr_IF_21 & ((\regs[0][0]~q )))))

	.dataa(Instr_IF_22),
	.datab(Instr_IF_21),
	.datac(\regs[1][0]~q ),
	.datad(\regs[0][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~634_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~634 .lut_mask = 16'hD9C8;
defparam \rfif.rdat1[0]~634 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \rfif.rdat1[0]~635 (
// Equation(s):
// \rfif.rdat1[0]~635_combout  = (Instr_IF_22 & ((\rfif.rdat1[0]~634_combout  & (\regs[3][0]~q )) # (!\rfif.rdat1[0]~634_combout  & ((\regs[2][0]~q ))))) # (!Instr_IF_22 & (((\rfif.rdat1[0]~634_combout ))))

	.dataa(Instr_IF_22),
	.datab(\regs[3][0]~q ),
	.datac(\regs[2][0]~q ),
	.datad(\rfif.rdat1[0]~634_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~635_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~635 .lut_mask = 16'hDDA0;
defparam \rfif.rdat1[0]~635 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N3
dffeas \regs[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[5][0] .is_wysiwyg = "true";
defparam \regs[5][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N15
dffeas \regs[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(input_a14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regs[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \regs[4][0] .is_wysiwyg = "true";
defparam \regs[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \rfif.rdat1[0]~632 (
// Equation(s):
// \rfif.rdat1[0]~632_combout  = (Instr_IF_21 & (Instr_IF_22)) # (!Instr_IF_21 & ((Instr_IF_22 & ((\regs[6][0]~q ))) # (!Instr_IF_22 & (\regs[4][0]~q ))))

	.dataa(Instr_IF_21),
	.datab(Instr_IF_22),
	.datac(\regs[4][0]~q ),
	.datad(\regs[6][0]~q ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~632_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~632 .lut_mask = 16'hDC98;
defparam \rfif.rdat1[0]~632 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \rfif.rdat1[0]~633 (
// Equation(s):
// \rfif.rdat1[0]~633_combout  = (Instr_IF_21 & ((\rfif.rdat1[0]~632_combout  & ((\regs[7][0]~q ))) # (!\rfif.rdat1[0]~632_combout  & (\regs[5][0]~q )))) # (!Instr_IF_21 & (((\rfif.rdat1[0]~632_combout ))))

	.dataa(Instr_IF_21),
	.datab(\regs[5][0]~q ),
	.datac(\regs[7][0]~q ),
	.datad(\rfif.rdat1[0]~632_combout ),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~633_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~633 .lut_mask = 16'hF588;
defparam \rfif.rdat1[0]~633 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \rfif.rdat1[0]~636 (
// Equation(s):
// \rfif.rdat1[0]~636_combout  = (Instr_IF_24 & (((Instr_IF_23)))) # (!Instr_IF_24 & ((Instr_IF_23 & ((\rfif.rdat1[0]~633_combout ))) # (!Instr_IF_23 & (\rfif.rdat1[0]~635_combout ))))

	.dataa(\rfif.rdat1[0]~635_combout ),
	.datab(Instr_IF_24),
	.datac(\rfif.rdat1[0]~633_combout ),
	.datad(Instr_IF_23),
	.cin(gnd),
	.combout(\rfif.rdat1[0]~636_combout ),
	.cout());
// synopsys translate_off
defparam \rfif.rdat1[0]~636 .lut_mask = 16'hFC22;
defparam \rfif.rdat1[0]~636 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	Memwrite_EX,
	MemToReg_EX,
	always0,
	devpor,
	devclrn,
	devoe);
input 	Memwrite_EX;
input 	MemToReg_EX;
output 	always0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// always0 = (MemToReg_EX1) # (Memwrite_EX1)

	.dataa(gnd),
	.datab(gnd),
	.datac(MemToReg_EX),
	.datad(Memwrite_EX),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hFFF0;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	\ramif.ramaddr ,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	ramWEN,
	ramREN,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr16,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	syiftbCTRL,
	syifaddr_25,
	syifaddr_24,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	ramWEN;
input 	ramREN;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr16;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	syiftbCTRL;
input 	syifaddr_25;
input 	syifaddr_24;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \Equal2~2_combout ;
wire \Equal2~5_combout ;
wire \Equal2~11_combout ;
wire \Equal2~15_combout ;
wire \Equal2~16_combout ;
wire \Equal2~17_combout ;
wire \always0~0_combout ;
wire \addr[8]~feeder_combout ;
wire \always0~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~3_combout ;
wire \Equal2~1_combout ;
wire \Equal2~4_combout ;
wire \Equal2~12_combout ;
wire \Equal2~13_combout ;
wire \Equal2~10_combout ;
wire \Equal2~14_combout ;
wire \Equal2~19_combout ;
wire \Equal2~18_combout ;
wire \Equal2~20_combout ;
wire \Equal2~21_combout ;
wire \Equal2~6_combout ;
wire \Equal2~8_combout ;
wire \Equal2~7_combout ;
wire \Equal2~9_combout ;
wire \Equal2~22_combout ;
wire [1:0] en;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3,ramaddr,ramaddr1}),
	.ramaddr(ramaddr12),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr16),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X60_Y32_N25
dffeas \addr[2] (
	.clk(CLK),
	.d(ramaddr1),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N13
dffeas \addr[4] (
	.clk(CLK),
	.d(ramaddr3),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N15
dffeas \addr[5] (
	.clk(CLK),
	.d(ramaddr2),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (addr[5] & (\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout )))) # (!addr[5] & (!\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout ))))

	.dataa(addr[5]),
	.datab(addr[4]),
	.datac(ramaddr2),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h8421;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \addr[6] (
	.clk(CLK),
	.d(ramaddr5),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N5
dffeas \addr[8] (
	.clk(CLK),
	.d(\addr[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N3
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr6),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (addr[8] & (\ramaddr~19_combout  & (addr[9] $ (!\ramaddr~17_combout )))) # (!addr[8] & (!\ramaddr~19_combout  & (addr[9] $ (!\ramaddr~17_combout ))))

	.dataa(addr[8]),
	.datab(ramaddr7),
	.datac(addr[9]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'h9009;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N9
dffeas \addr[10] (
	.clk(CLK),
	.d(ramaddr9),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N15
dffeas \addr[13] (
	.clk(CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N11
dffeas \addr[14] (
	.clk(CLK),
	.d(ramaddr13),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N25
dffeas \addr[16] (
	.clk(CLK),
	.d(\ramif.ramaddr [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N29
dffeas \addr[18] (
	.clk(CLK),
	.d(\ramif.ramaddr [18]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N23
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \Equal2~11 (
// Equation(s):
// \Equal2~11_combout  = (addr[18] & (\ramaddr~39_combout  & (addr[19] $ (!\ramaddr~37_combout )))) # (!addr[18] & (!\ramaddr~39_combout  & (addr[19] $ (!\ramaddr~37_combout ))))

	.dataa(addr[18]),
	.datab(addr[19]),
	.datac(\ramif.ramaddr [19]),
	.datad(\ramif.ramaddr [18]),
	.cin(gnd),
	.combout(\Equal2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~11 .lut_mask = 16'h8241;
defparam \Equal2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N19
dffeas \addr[20] (
	.clk(CLK),
	.d(\ramif.ramaddr [20]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N29
dffeas \addr[22] (
	.clk(CLK),
	.d(\ramif.ramaddr [22]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \addr[25] (
	.clk(CLK),
	.d(\ramif.ramaddr [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \Equal2~15 (
// Equation(s):
// \Equal2~15_combout  = addr[25] $ (((\syif.tbCTRL~input_o  & \syif.addr[25]~input_o )))

	.dataa(syiftbCTRL),
	.datab(gnd),
	.datac(addr[25]),
	.datad(syifaddr_25),
	.cin(gnd),
	.combout(\Equal2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~15 .lut_mask = 16'h5AF0;
defparam \Equal2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N13
dffeas \addr[24] (
	.clk(CLK),
	.d(\ramif.ramaddr [24]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \Equal2~16 (
// Equation(s):
// \Equal2~16_combout  = addr[24] $ (((\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~49_combout )))))

	.dataa(addr[24]),
	.datab(syifaddr_24),
	.datac(syiftbCTRL),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\Equal2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~16 .lut_mask = 16'h656A;
defparam \Equal2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \Equal2~17 (
// Equation(s):
// \Equal2~17_combout  = (!\Equal2~16_combout  & (\Equal2~15_combout  $ (((\syif.tbCTRL~input_o ) # (!\ramaddr~48_combout )))))

	.dataa(ramaddr14),
	.datab(syiftbCTRL),
	.datac(\Equal2~15_combout ),
	.datad(\Equal2~16_combout ),
	.cin(gnd),
	.combout(\Equal2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~17 .lut_mask = 16'h002D;
defparam \Equal2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N9
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N27
dffeas \addr[30] (
	.clk(CLK),
	.d(\ramif.ramaddr [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N27
dffeas \en[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramREN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N7
dffeas \en[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramWEN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (en[0] & ((\ramREN~0_combout  $ (en[1])) # (!\ramWEN~0_combout ))) # (!en[0] & ((\ramWEN~0_combout ) # (\ramREN~0_combout  $ (en[1]))))

	.dataa(en[0]),
	.datab(ramREN),
	.datac(en[1]),
	.datad(ramWEN),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h7DBE;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \addr[8]~feeder (
// Equation(s):
// \addr[8]~feeder_combout  = \ramaddr~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr7),
	.cin(gnd),
	.combout(\addr[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[8]~feeder .lut_mask = 16'hFF00;
defparam \addr[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((\Equal2~22_combout  & ((!\ramREN~0_combout ) # (!\ramWEN~0_combout )))) # (!\nRST~input_o )

	.dataa(ramWEN),
	.datab(nRST),
	.datac(ramREN),
	.datad(\Equal2~22_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h7F33;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & (ram_block3a331)) # (!address_reg_a_0 & ((ram_block3a110)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'h8A80;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hD800;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N18
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & ((ram_block3a351))) # (!address_reg_a_0 & (ram_block3a310))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'hE400;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N20
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hFD75;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N18
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hE020;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N4
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & ((ram_block3a381))) # (!address_reg_a_0 & (ram_block3a64))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & ((ram_block3a391))) # (!address_reg_a_0 & (ram_block3a71))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hFB3B;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & ((ram_block3a401))) # (!address_reg_a_0 & (ram_block3a81))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hC840;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N8
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & (ram_block3a421)) # (!address_reg_a_0 & ((ram_block3a101)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hB800;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & ((ram_block3a431))) # (!address_reg_a_0 & (ram_block3a112))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hEF2F;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & (ram_block3a441)) # (!address_reg_a_0 & ((ram_block3a121)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hB8FF;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hFD75;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & ((ram_block3a461))) # (!address_reg_a_0 & (ram_block3a141))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'hC808;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & (ram_block3a471)) # (!address_reg_a_0 & ((ram_block3a151)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hDFD5;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & ((ram_block3a481))) # (!address_reg_a_0 & (ram_block3a161))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \ramif.ramload[17]~17 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & ((ram_block3a491))) # (!address_reg_a_0 & (ram_block3a171))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~17 .lut_mask = 16'hA808;
defparam \ramif.ramload[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \ramif.ramload[18]~18 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & (ram_block3a501)) # (!address_reg_a_0 & ((ram_block3a181)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~18 .lut_mask = 16'hB800;
defparam \ramif.ramload[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \ramif.ramload[19]~19 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & ((ram_block3a512))) # (!address_reg_a_0 & (ram_block3a191))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~19 .lut_mask = 16'hA808;
defparam \ramif.ramload[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N8
cycloneive_lcell_comb \ramif.ramload[20]~20 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & (ram_block3a521)) # (!address_reg_a_0 & ((ram_block3a201)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~20 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \ramif.ramload[21]~21 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & (ram_block3a531)) # (!address_reg_a_0 & ((ram_block3a212)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~21 .lut_mask = 16'hD080;
defparam \ramif.ramload[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \ramif.ramload[22]~22 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~22 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \ramif.ramload[23]~23 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & ((ram_block3a551))) # (!address_reg_a_0 & (ram_block3a231))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~23 .lut_mask = 16'hFD75;
defparam \ramif.ramload[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \ramif.ramload[24]~24 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~24 .lut_mask = 16'hA088;
defparam \ramif.ramload[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \ramif.ramload[25]~25 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & (ram_block3a571)) # (!address_reg_a_0 & ((ram_block3a251)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~25 .lut_mask = 16'hDFD5;
defparam \ramif.ramload[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \ramif.ramload[26]~26 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & (ram_block3a581)) # (!address_reg_a_0 & ((ram_block3a261)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~26 .lut_mask = 16'hA280;
defparam \ramif.ramload[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \ramif.ramload[27]~27 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~27 .lut_mask = 16'hBFB3;
defparam \ramif.ramload[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \ramif.ramload[28]~28 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & ((ram_block3a601))) # (!address_reg_a_0 & (ram_block3a281))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~28 .lut_mask = 16'hFD75;
defparam \ramif.ramload[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \ramif.ramload[29]~29 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~29 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \ramif.ramload[30]~30 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & ((ram_block3a621))) # (!address_reg_a_0 & (ram_block3a301))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~30 .lut_mask = 16'hC840;
defparam \ramif.ramload[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \ramif.ramload[31]~31 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~31 .lut_mask = 16'hFD75;
defparam \ramif.ramload[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\always0~0_combout ) # (((\ramREN~0_combout  & \ramWEN~0_combout )) # (!\Equal2~22_combout ))

	.dataa(\always0~0_combout ),
	.datab(ramREN),
	.datac(ramWEN),
	.datad(\Equal2~22_combout ),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'hEAFF;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N23
dffeas \addr[1] (
	.clk(CLK),
	.d(\ramif.ramaddr [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N21
dffeas \addr[0] (
	.clk(CLK),
	.d(\ramif.ramaddr [0]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (\ramaddr~1_combout  & (addr[1] & (addr[0] $ (!\ramaddr~3_combout )))) # (!\ramaddr~1_combout  & (!addr[1] & (addr[0] $ (!\ramaddr~3_combout ))))

	.dataa(\ramif.ramaddr [1]),
	.datab(addr[1]),
	.datac(addr[0]),
	.datad(\ramif.ramaddr [0]),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h9009;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N5
dffeas \addr[7] (
	.clk(CLK),
	.d(ramaddr4),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = (addr[6] & (\ramaddr~15_combout  & (addr[7] $ (!\ramaddr~13_combout )))) # (!addr[6] & (!\ramaddr~15_combout  & (addr[7] $ (!\ramaddr~13_combout ))))

	.dataa(addr[6]),
	.datab(addr[7]),
	.datac(ramaddr4),
	.datad(ramaddr5),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h8241;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N15
dffeas \addr[3] (
	.clk(CLK),
	.d(ramaddr),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (addr[2] & (\ramaddr~7_combout  & (addr[3] $ (!\ramaddr~5_combout )))) # (!addr[2] & (!\ramaddr~7_combout  & (addr[3] $ (!\ramaddr~5_combout ))))

	.dataa(addr[2]),
	.datab(addr[3]),
	.datac(ramaddr),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h8241;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// \Equal2~4_combout  = (\Equal2~2_combout  & (\Equal2~0_combout  & (\Equal2~3_combout  & \Equal2~1_combout )))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~0_combout ),
	.datac(\Equal2~3_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'h8000;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N13
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \Equal2~12 (
// Equation(s):
// \Equal2~12_combout  = (addr[20] & (\ramaddr~43_combout  & (addr[21] $ (!\ramaddr~41_combout )))) # (!addr[20] & (!\ramaddr~43_combout  & (addr[21] $ (!\ramaddr~41_combout ))))

	.dataa(addr[20]),
	.datab(\ramif.ramaddr [20]),
	.datac(addr[21]),
	.datad(\ramif.ramaddr [21]),
	.cin(gnd),
	.combout(\Equal2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~12 .lut_mask = 16'h9009;
defparam \Equal2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N31
dffeas \addr[23] (
	.clk(CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \Equal2~13 (
// Equation(s):
// \Equal2~13_combout  = (addr[22] & (\ramaddr~47_combout  & (addr[23] $ (!\ramaddr~45_combout )))) # (!addr[22] & (!\ramaddr~47_combout  & (addr[23] $ (!\ramaddr~45_combout ))))

	.dataa(addr[22]),
	.datab(addr[23]),
	.datac(\ramif.ramaddr [23]),
	.datad(\ramif.ramaddr [22]),
	.cin(gnd),
	.combout(\Equal2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~13 .lut_mask = 16'h8241;
defparam \Equal2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N31
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \Equal2~10 (
// Equation(s):
// \Equal2~10_combout  = (addr[16] & (\ramaddr~35_combout  & (addr[17] $ (!\ramaddr~33_combout )))) # (!addr[16] & (!\ramaddr~35_combout  & (addr[17] $ (!\ramaddr~33_combout ))))

	.dataa(addr[16]),
	.datab(addr[17]),
	.datac(\ramif.ramaddr [17]),
	.datad(\ramif.ramaddr [16]),
	.cin(gnd),
	.combout(\Equal2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~10 .lut_mask = 16'h8241;
defparam \Equal2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \Equal2~14 (
// Equation(s):
// \Equal2~14_combout  = (\Equal2~11_combout  & (\Equal2~12_combout  & (\Equal2~13_combout  & \Equal2~10_combout )))

	.dataa(\Equal2~11_combout ),
	.datab(\Equal2~12_combout ),
	.datac(\Equal2~13_combout ),
	.datad(\Equal2~10_combout ),
	.cin(gnd),
	.combout(\Equal2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~14 .lut_mask = 16'h8000;
defparam \Equal2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N23
dffeas \addr[28] (
	.clk(CLK),
	.d(\ramif.ramaddr [28]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \Equal2~19 (
// Equation(s):
// \Equal2~19_combout  = (addr[29] & (\ramaddr~55_combout  & (addr[28] $ (!\ramaddr~57_combout )))) # (!addr[29] & (!\ramaddr~55_combout  & (addr[28] $ (!\ramaddr~57_combout ))))

	.dataa(addr[29]),
	.datab(addr[28]),
	.datac(\ramif.ramaddr [29]),
	.datad(\ramif.ramaddr [28]),
	.cin(gnd),
	.combout(\Equal2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~19 .lut_mask = 16'h8421;
defparam \Equal2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N3
dffeas \addr[26] (
	.clk(CLK),
	.d(\ramif.ramaddr [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \Equal2~18 (
// Equation(s):
// \Equal2~18_combout  = (addr[27] & (\ramaddr~51_combout  & (\ramaddr~53_combout  $ (!addr[26])))) # (!addr[27] & (!\ramaddr~51_combout  & (\ramaddr~53_combout  $ (!addr[26]))))

	.dataa(addr[27]),
	.datab(\ramif.ramaddr [26]),
	.datac(addr[26]),
	.datad(\ramif.ramaddr [27]),
	.cin(gnd),
	.combout(\Equal2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~18 .lut_mask = 16'h8241;
defparam \Equal2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \Equal2~20 (
// Equation(s):
// \Equal2~20_combout  = (addr[30] & (\ramaddr~61_combout  & (addr[31] $ (!\ramaddr~59_combout )))) # (!addr[30] & (!\ramaddr~61_combout  & (addr[31] $ (!\ramaddr~59_combout ))))

	.dataa(addr[30]),
	.datab(addr[31]),
	.datac(\ramif.ramaddr [31]),
	.datad(\ramif.ramaddr [30]),
	.cin(gnd),
	.combout(\Equal2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~20 .lut_mask = 16'h8241;
defparam \Equal2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \Equal2~21 (
// Equation(s):
// \Equal2~21_combout  = (\Equal2~17_combout  & (\Equal2~19_combout  & (\Equal2~18_combout  & \Equal2~20_combout )))

	.dataa(\Equal2~17_combout ),
	.datab(\Equal2~19_combout ),
	.datac(\Equal2~18_combout ),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\Equal2~21_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~21 .lut_mask = 16'h8000;
defparam \Equal2~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N3
dffeas \addr[11] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (addr[10] & (\ramaddr~23_combout  & (addr[11] $ (!\ramaddr~21_combout )))) # (!addr[10] & (!\ramaddr~23_combout  & (addr[11] $ (!\ramaddr~21_combout ))))

	.dataa(addr[10]),
	.datab(addr[11]),
	.datac(ramaddr9),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h8421;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y29_N29
dffeas \addr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N28
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// \Equal2~8_combout  = (addr[14] & (\ramaddr~31_combout  & (\ramaddr~29_combout  $ (addr[15])))) # (!addr[14] & (!\ramaddr~31_combout  & (\ramaddr~29_combout  $ (addr[15]))))

	.dataa(addr[14]),
	.datab(ramaddr12),
	.datac(addr[15]),
	.datad(ramaddr13),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h2814;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y29_N13
dffeas \addr[12] (
	.clk(CLK),
	.d(ramaddr11),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N16
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// \Equal2~7_combout  = (addr[13] & (\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout )))) # (!addr[13] & (!\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout ))))

	.dataa(addr[13]),
	.datab(addr[12]),
	.datac(ramaddr10),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'h8421;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// \Equal2~9_combout  = (\Equal2~5_combout  & (\Equal2~6_combout  & (\Equal2~8_combout  & \Equal2~7_combout )))

	.dataa(\Equal2~5_combout ),
	.datab(\Equal2~6_combout ),
	.datac(\Equal2~8_combout ),
	.datad(\Equal2~7_combout ),
	.cin(gnd),
	.combout(\Equal2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h8000;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Equal2~22 (
// Equation(s):
// \Equal2~22_combout  = (\Equal2~4_combout  & (\Equal2~14_combout  & (\Equal2~21_combout  & \Equal2~9_combout )))

	.dataa(\Equal2~4_combout ),
	.datab(\Equal2~14_combout ),
	.datac(\Equal2~21_combout ),
	.datad(\Equal2~9_combout ),
	.cin(gnd),
	.combout(\Equal2~22_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~22 .lut_mask = 16'h8000;
defparam \Equal2~22 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_a[0]~feeder_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X15_Y30_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001802C7EA14A7EF95C00000000000000000000000000000A242111E008528F7260;
// synopsys translate_on

// Location: M9K_X37_Y40_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y41_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D4AE6429116B3C8A000000000000000000000000000012242108900D12808390;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000961CA470728D97800000000000000000000000000000172E7BD1C323272F6867;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009F20E64C2468E52000000000000000000000000000022346308C62632A08083;
// synopsys translate_on

// Location: M9K_X37_Y28_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y27_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060B81842D24565BE000000000000000000000000000002242101022202208083;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000056414512D6B00448000000000000000000000000000002246308006652AF7263;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001003088D801A0F827000000000000000000000000000012042100402202200113;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220A200403;
// synopsys translate_on

// Location: M9K_X37_Y29_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220230080F;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y30_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002202300003;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210800265A2A2233;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022C2043;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022F5213;
// synopsys translate_on

// Location: M9K_X78_Y29_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y28_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000224A200503;
// synopsys translate_on

// Location: M9K_X78_Y40_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y39_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002242206063;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000205A122003613254042;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006C0340C001602060001;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060C3180001703286867;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C38C6E09B6D7701203;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y27_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A0832F000B;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002A142119BCBBAB600000;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y41_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E403004A40002000000;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E5CB187BC004B601000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021830C680DB793600400;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000CB783600310;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X15_Y31_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007CFBDE639B287F0888F;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010E1C6264AD282C08088;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008100011B00926100807;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X15_Y34_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078F3DE001B007700807;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X15_Y33_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000C18426089282400008;
// synopsys translate_on

// Location: FF_X59_Y28_N25
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(\address_reg_a[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N13
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N24
cycloneive_lcell_comb \address_reg_a[0]~feeder (
// Equation(s):
// \address_reg_a[0]~feeder_combout  = \ramaddr~29_wirecell_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\address_reg_a[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_a[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_a[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (always1 & (!\ramaddr~29_combout  & !\ramWEN~0_combout ))

	.dataa(always1),
	.datab(ramaddr),
	.datac(ramWEN),
	.datad(gnd),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0202;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(ramaddr),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h4040;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X67_Y36_N22
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (ram_rom_addr_reg_13 & sdr)))

	.dataa(irf_reg_2_1),
	.datab(state_5),
	.datac(ram_rom_addr_reg_13),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N16
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (!ram_rom_addr_reg_13 & sdr)))

	.dataa(irf_reg_2_1),
	.datab(state_5),
	.datac(ram_rom_addr_reg_13),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h0800;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~2_combout ;
wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \Add1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[26]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[2]~42_combout ;
wire \ram_rom_addr_reg[2]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X68_Y36_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X68_Y36_N27
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~6_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h8F0F;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N29
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N17
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N31
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N5
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N7
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N9
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N11
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N13
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N15
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N17
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N19
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N21
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N23
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N25
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N27
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N29
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[2]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N23
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N13
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N15
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N29
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N3
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N5
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N31
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N21
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N27
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y33_N9
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N29
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N27
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N25
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N11
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N5
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N23
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N21
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N31
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N9
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N15
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N21
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N23
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N31
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N27
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N9
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N15
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N5
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N3
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N25
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N19
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N29
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[26]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N13
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_0),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N27
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N1
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N31
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N10
cycloneive_lcell_comb \tdo~1 (
	.dataa(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(\tdo~0_combout ),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hAFA0;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N12
cycloneive_lcell_comb \sdr~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(node_ena_1),
	.datad(gnd),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h5050;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N28
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N16
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a0),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a32),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_2_1),
	.datab(state_4),
	.datac(sdr),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC080;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Add1~2_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h08B8;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N5
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h33CC;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h070F;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N3
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N1
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~8_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N29
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~10_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N31
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N8
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[2]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N6
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Equal1~0_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hF000;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N26
cycloneive_lcell_comb \process_0~2 (
	.dataa(\Equal1~1_combout ),
	.datab(ir_in[3]),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h1333;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \ram_rom_data_reg[26]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\process_0~2_combout ),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~32 .lut_mask = 16'hFF0F;
defparam \ram_rom_data_reg[26]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(ram_rom_addr_reg_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(ram_rom_addr_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h5A5A;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N18
cycloneive_lcell_comb \process_0~3 (
	.dataa(virtual_ir_scan_reg),
	.datab(ir_in[3]),
	.datac(node_ena_1),
	.datad(state_4),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h4000;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N24
cycloneive_lcell_comb \ram_rom_addr_reg[2]~42 (
	.dataa(\Equal1~1_combout ),
	.datab(\process_0~3_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[2]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~42 .lut_mask = 16'hCECC;
defparam \ram_rom_addr_reg[2]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N30
cycloneive_lcell_comb \ram_rom_addr_reg[2]~43 (
	.dataa(irf_reg_2_1),
	.datab(\ram_rom_addr_reg[2]~42_combout ),
	.datac(state_8),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[2]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~43 .lut_mask = 16'hECCC;
defparam \ram_rom_addr_reg[2]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a1),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a33),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a2),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a34),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a3),
	.datab(ram_block3a35),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a4),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a36),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N2
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a5),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a37),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N4
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a6),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a38),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a39),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a7),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N20
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a8),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a40),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a9),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a41),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a42),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a10),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(ram_block3a43),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a11),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(ram_block3a44),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a12),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a13),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a45),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(ram_block3a14),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a46),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a15),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a47),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(ram_block3a48),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a16),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a17),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a49),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(ram_block3a50),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a18),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a51),
	.datac(gnd),
	.datad(ram_block3a19),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a52),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a20),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a21),
	.datac(gnd),
	.datad(ram_block3a53),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a54),
	.datac(gnd),
	.datad(ram_block3a22),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(ram_block3a55),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(ram_block3a24),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a25),
	.datab(ram_block3a57),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a58),
	.datab(ram_block3a26),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a59),
	.datac(gnd),
	.datad(ram_block3a27),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a28),
	.datab(ram_block3a60),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a29),
	.datac(gnd),
	.datad(ram_block3a61),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a30),
	.datab(ram_block3a62),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(ram_block3a63),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N14
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFFF0;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N0
cycloneive_lcell_comb \process_0~1 (
	.dataa(virtual_ir_scan_reg),
	.datab(node_ena_1),
	.datac(state_5),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h4000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N26
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N30
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N2
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(gnd),
	.datab(node_ena_1),
	.datac(\bypass_reg_out~q ),
	.datad(altera_internal_jtag),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hFC30;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N3
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N20
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(\bypass_reg_out~q ),
	.datac(ram_rom_data_reg_0),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hF0E4;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \word_counter[1]~9_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \word_counter[3]~13_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[3]~19_combout ;
wire \word_counter[3]~14_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \word_counter[3]~15_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[2]~6_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: FF_X67_Y38_N23
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[3]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[3]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N22
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(word_counter[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h5A5F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hAB08;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N4
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(state_4),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h000B;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N6
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(gnd),
	.datab(\WORD_SR~7_combout ),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h000C;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N10
cycloneive_lcell_comb \word_counter[3]~13 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[1]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\word_counter[3]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[3]~13 .lut_mask = 16'hFBFF;
defparam \word_counter[3]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N10
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hF784;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N0
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(\WORD_SR~10_combout ),
	.datab(gnd),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hA5A0;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N13
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N8
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(virtual_ir_scan_reg),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hC0C0;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N20
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N14
cycloneive_lcell_comb \word_counter[3]~19 (
	.dataa(\word_counter[3]~13_combout ),
	.datab(virtual_ir_scan_reg),
	.datac(state_8),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\word_counter[3]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[3]~19 .lut_mask = 16'hC0D5;
defparam \word_counter[3]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N0
cycloneive_lcell_comb \word_counter[3]~14 (
	.dataa(state_3),
	.datab(\clear_signal~combout ),
	.datac(state_4),
	.datad(sdr),
	.cin(gnd),
	.combout(\word_counter[3]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[3]~14 .lut_mask = 16'hCECC;
defparam \word_counter[3]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N21
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[3]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[3]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N24
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X67_Y38_N25
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[3]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[3]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N26
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N28
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(gnd),
	.datab(word_counter[4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hC3C3;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X67_Y38_N29
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[3]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[3]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N27
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[3]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[3]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N18
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h2000;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(altera_internal_jtag),
	.datab(\WORD_SR~13_combout ),
	.datac(word_counter[0]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hAA0C;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N18
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(gnd),
	.datab(virtual_ir_scan_reg),
	.datac(state_8),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h3F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N2
cycloneive_lcell_comb \WORD_SR[2]~6 (
	.dataa(state_3),
	.datab(\clear_signal~combout ),
	.datac(state_4),
	.datad(sdr),
	.cin(gnd),
	.combout(\WORD_SR[2]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[2]~6 .lut_mask = 16'hFECC;
defparam \WORD_SR[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N19
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N16
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(\WORD_SR~11_combout ),
	.datab(state_4),
	.datac(\clear_signal~combout ),
	.datad(WORD_SR[3]),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h0E02;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N17
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N30
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(state_4),
	.datac(\clear_signal~combout ),
	.datad(WORD_SR[2]),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h0E0A;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N31
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N12
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h3005;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~3_combout ),
	.datab(gnd),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hAAA0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N12
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(state_4),
	.datac(\clear_signal~combout ),
	.datad(\WORD_SR~4_combout ),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h0B08;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
