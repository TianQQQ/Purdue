/*
  Eric Villasenor
  evillase@gmail.com

  this block is the coherence protocol
  and artibtration for ram
*/

// interface include
`include "control_unit_if.vh"

// memory types
`include "cpu_types_pkg.vh"
 import cpu_types_pkg::*;

module control_unit (
  control_unit_if cuif
);


	/***************************************************************
	---------------------<Pseudo Instructions>-----------------------
	PUSH   $rs           $29 <= $29 - 4; Mem[$29+0] <= R[rs] (sub+sw)
	POP    $rt           R[rt] <= Mem[$29+0]; $29 <= $29 + 4 (add+lw)
	NOP                  Nop
	-----------------------------------------------------------------
	-----------------------------------------------------------------
	org  Addr         Set the base address for the code to follow 
	chw  #            Assign value to half word memory
	cfw  #            Assign value to word of memory
	**************************************************************/


   always_comb
     begin
	cuif.jump = 3'b000; cuif.RegDst = 2'b00; cuif.RegWen = 0; cuif.ALUSrc = 3'b000; cuif.ALUOP = ALU_SLL;cuif.MemToReg = 0; cuif.PcToReg = 0;cuif.MemWrite = 0; cuif.careOF = 0;cuif.halt = 0;

	cuif.input_hazard_Reg_ID = 0;

	unique casez(cuif.Instr[31:26])

		/****************************************************************
		---------------------<R-type Instructions>-----------------------
		ADDU   $rd,$rs,$rt   R[rd] <= R[rs] + R[rt] (unchecked overflow)
		ADD    $rd,$rs,$rt   R[rd] <= R[rs] + R[rt]
		AND    $rd,$rs,$rt   R[rd] <= R[rs] AND R[rt]
		JR     $rs           PC <= R[rs]
		NOR    $rd,$rs,$rt   R[rd] <= ~(R[rs] OR R[rt])
		OR     $rd,$rs,$rt   R[rd] <= R[rs] OR R[rt]
		SLT    $rd,$rs,$rt   R[rd] <= (R[rs] < R[rt]) ? 1 : 0
		SLTU   $rd,$rs,$rt   R[rd] <= (R[rs] < R[rt]) ? 1 : 0
		SLL    $rd,$rs,shamt R[rd] <= R[rs] << shamt
		SRL    $rd,$rs,shamt R[rd] <= R[rs] >> shamt
		SUBU   $rd,$rs,$rt   R[rd] <= R[rs] - R[rt] (unchecked overflow)
		SUB    $rd,$rs,$rt   R[rd] <= R[rs] - R[rt]
		XOR    $rd,$rs,$rt   R[rd] <= R[rs] XOR R[rt]
		*****************************************************************/

	  RTYPE: //r instructions
	    begin
	       cuif.input_hazard_Reg_ID = 1;

	       unique casez(cuif.Instr[5:0])
		 SLL:
		   begin
		      cuif.ALUOP = ALU_SLL;
		      cuif.ALUSrc = 3'b100;
		      cuif.RegWen = 1;
		   end

		 SRL:
		   begin
		      cuif.ALUOP = ALU_SRL;
		      cuif.ALUSrc = 3'b100;
		      cuif.RegWen = 1;
		   end

		 JR:
		   begin
		      cuif.jump = 3'b010;
		   end

		 ADD:
		   begin
		      cuif.ALUOP = ALU_ADD;
		      cuif.RegWen = 1;
		      cuif.careOF = 1;
		   end

		 SUB:
		   begin
		      cuif.ALUOP = ALU_SUB;
		      cuif.RegWen = 1;
		      cuif.careOF = 1;
		   end

		 SUBU:
		   begin
		      cuif.ALUOP = ALU_SUB;
		      cuif.RegWen = 1;
		   end

		 AND:
		   begin
		      cuif.ALUOP = ALU_AND;
		      cuif.RegWen = 1;
		   end

		 OR:
		   begin
		      cuif.ALUOP = ALU_OR;
		      cuif.RegWen = 1;
		   end

		 XOR:
		   begin
		      cuif.ALUOP = ALU_XOR;
		      cuif.RegWen = 1;
		   end

		 NOR:
		   begin
		      cuif.ALUOP = ALU_NOR;
		      cuif.RegWen = 1;
		   end

		 SLT:
		   begin
		      cuif.ALUOP = ALU_SLT;
		      cuif.RegWen = 1;
		   end
 		 ADDU:
		   begin
		      cuif.ALUOP = ALU_ADD;
		      cuif.RegWen = 1;
		   end
		 SLTU:
		   begin
		      cuif.ALUOP = ALU_SLTU;
		      cuif.RegWen = 1;
		   end

	       endcase
	    end




	/****************************************************************************************
	---------------------<I-type Instructions>-----------------------
	ADDIU  $rt,$rs,imm   R[rt] <= R[rs] + SignExtImm (unchecked overflow)
	ADDI   $rt,$rs,imm   R[rt] <= R[rs] + SignExtImm
	ANDI   $rt,$rs,imm   R[rt] <= R[rs] & ZeroExtImm
	BEQ    $rs,$rt,label PC <= (R[rs] == R[rt]) ? npc+BranchAddr : npc
	BNE    $rs,$rt,label PC <= (R[rs] != R[rt]) ? npc+BranchAddr : npc
	LUI    $rt,imm       R[rt] <= {imm,16b'0}
	LW     $rt,imm($rs)  R[rt] <= M[R[rs] + SignExtImm]
	ORI    $rt,$rs,imm   R[rt] <= R[rs] OR ZeroExtImm
	SLTI   $rt,$rs,imm   R[rt] <= (R[rs] < SignExtImm) ? 1 : 0
	SLTIU  $rt,$rs,imm   R[rt] <= (R[rs] < SignExtImm) ? 1 : 0
	SW     $rt,imm($rs)  M[R[rs] + SignExtImm] <= R[rt]
	LL     $rt,imm($rs)  R[rt] <= M[R[rs] + SignExtImm]; rmwstate <= addr
	SC     $rt,imm($rs)  if (rmw) M[R[rs] + SignExtImm] <= R[rt], R[rt] <= 1 else R[rt] <= 0
	XORI   $rt,$rs,imm   R[rt] <= R[rs] XOR ZeroExtImm
	****************************************************************************************/
	  //itype
	  BEQ:
	    begin
	       cuif.jump = 3'b011;
	       cuif.ALUOP = ALU_SUB;
	    end

	  BNE:
	    begin
	       cuif.jump = 3'b100;
	       cuif.ALUOP = ALU_SUB;
	    end

	  ADDI:
	    begin
	       cuif.ALUOP = ALU_ADD;
	       cuif.ALUSrc = 3'b001;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	       cuif.careOF = 1;
	    end

	  ADDIU:
	    begin
	       cuif.ALUOP = ALU_ADD;
	       cuif.ALUSrc = 3'b001;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  SLTI:
	    begin
	       cuif.ALUOP = ALU_SLT;
	       cuif.ALUSrc = 3'b001;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  SLTIU:
	    begin
	       cuif.ALUOP = ALU_SLTU;
	       cuif.ALUSrc = 3'b001;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end


	  SW:
	    begin
	       cuif.ALUOP = ALU_ADD;
	       cuif.ALUSrc = 3'b001;
	       cuif.MemWrite = 1;
	       cuif.input_hazard_Reg_ID = 1;
	    end


	  ANDI:
	    begin
	       cuif.ALUOP = ALU_AND;
	       cuif.ALUSrc = 3'b010;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  ORI:
	    begin
	       cuif.ALUOP = ALU_OR;
	       cuif.ALUSrc = 3'b010;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  XORI:
	    begin
	       cuif.ALUOP = ALU_XOR;
	       cuif.ALUSrc = 3'b010;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  LUI:
	    begin
	       cuif.ALUOP = ALU_OR;
	       cuif.ALUSrc = 3'b011;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	    end

	  LW:
	    begin
	       cuif.ALUOP = ALU_ADD;
	       cuif.ALUSrc = 3'b001;
	       cuif.RegWen = 1;
	       cuif.RegDst = 2'b01;
	       cuif.MemToReg = 1;
	    end
	  


	/*******************************************************************
	---------------------<J-type Instructions>-----------------------
	J      label         PC <= JumpAddr
	JAL    label         R[31] <= npc; PC <= JumpAddr
	********************************************************************/
 


	  J:
	    begin
	       cuif.jump = 3'b001;
	    end

	  JAL:
	    begin
	       cuif.jump = 3'b001;
	       cuif.RegWen = 1'b1;
	       cuif.RegDst = 2'b10;
	       cuif.PcToReg = 1;
	    end


	/*---------------------<Other Instructions>------------------------
	HALT
	------------------------------------------------------------------*/
	  HALT:
	    begin
	       cuif.halt = 1;
	    end



	endcase
     end

endmodule
