/home/ecegrid/a/mg121/ece337/Lab2/source/adder_8bit.sv